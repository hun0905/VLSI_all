************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: part1_4
* View Name:     schematic
* Netlisted on:  Oct 30 23:18:57 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    part1_4
* View Name:    schematic
************************************************************************

.SUBCKT part1_4 A B C OUT VDD VSS
*.PININFO A:I B:I C:I OUT:O VDD:B VSS:B
MM5 OUT C VSS VSS NM W=1.5u L=180.00n
MM4 net5 B VSS VSS NM W=1.5u L=180.00n
MM3 OUT A net5 VSS NM W=1.5u L=180.00n
MM2 OUT C net21 VDD PM W=500.0n L=180.00n
MM1 net21 B VDD VDD PM W=500.0n L=180.00n
MM0 net21 A VDD VDD PM W=500.0n L=180.00n
.ENDS

