************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: nand4
* View Name:     schematic
* Netlisted on:  Jan 12 15:57:07 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    nand4
* View Name:    schematic
************************************************************************

.SUBCKT nand4 A B C D OUT VDD VSS
*.PININFO A:I B:I C:I D:I OUT:O VDD:B VSS:B
MM11 net030 D VSS VSS N_18 W=500.0n L=180.00n m=1
MM6 net40 C net030 VSS N_18 W=500.0n L=180.00n m=1
MM5 net44 B net40 VSS N_18 W=500.0n L=180.00n m=1
MM4 OUT A net44 VSS N_18 W=500.0n L=180.00n m=1
MM12 OUT D VDD VDD P_18 W=500.0n L=180.00n m=3
MM10 OUT A VDD VDD P_18 W=500.0n L=180.00n m=3
MM2 OUT C VDD VDD P_18 W=500.0n L=180.00n m=3
MM0 OUT B VDD VDD P_18 W=500.0n L=180.00n m=3
.ENDS

