* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT final_mux BL<1> BL<3> BL<5> BL<7> BL<0> BL<2> BL<4> BL<6> VSS VDD
** N=27 EP=10 IP=0 FDC=32
M0 15 1 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=5951 $Y=-13910 $D=0
M1 16 2 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=5951 $Y=-4410 $D=0
M2 BL<1> 1 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=6136 $Y=-15876 $D=0
M3 BL<0> 2 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=6136 $Y=-6376 $D=0
M4 18 3 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=8101 $Y=-13910 $D=0
M5 19 4 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=8101 $Y=-4410 $D=0
M6 BL<3> 3 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=8286 $Y=-15876 $D=0
M7 BL<2> 4 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=8286 $Y=-6376 $D=0
M8 21 5 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10251 $Y=-13910 $D=0
M9 22 6 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10251 $Y=-4410 $D=0
M10 BL<5> 5 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10436 $Y=-15876 $D=0
M11 BL<4> 6 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10436 $Y=-6376 $D=0
M12 24 7 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=12401 $Y=-13910 $D=0
M13 25 8 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=12401 $Y=-4410 $D=0
M14 BL<7> 7 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=12586 $Y=-15876 $D=0
M15 BL<6> 8 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=12586 $Y=-6376 $D=0
M16 15 1 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=5951 $Y=-12205 $D=1
M17 10 15 BL<1> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=5951 $Y=-9410 $D=1
M18 16 2 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=5951 $Y=-2705 $D=1
M19 10 16 BL<0> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=5951 $Y=90 $D=1
M20 18 3 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=8101 $Y=-12205 $D=1
M21 10 18 BL<3> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=8101 $Y=-9410 $D=1
M22 19 4 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=8101 $Y=-2705 $D=1
M23 10 19 BL<2> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=8101 $Y=90 $D=1
M24 21 5 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=10251 $Y=-12205 $D=1
M25 10 21 BL<5> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=10251 $Y=-9410 $D=1
M26 22 6 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=10251 $Y=-2705 $D=1
M27 10 22 BL<4> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=10251 $Y=90 $D=1
M28 24 7 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=12401 $Y=-12205 $D=1
M29 10 24 BL<7> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=12401 $Y=-9410 $D=1
M30 25 8 VDD VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=12401 $Y=-2705 $D=1
M31 10 25 BL<6> VDD P_18 L=1.8e-07 W=1.39e-06 AD=7.1145e-13 AS=7.1145e-13 PD=2.415e-06 PS=2.415e-06 $X=12401 $Y=90 $D=1
.ENDS
***************************************
