* File: hw2_part2_1_smaller.pex.spi
* Created: Fri Nov 12 00:13:50 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw2_part2_1_smaller.pex.spi.pex"
.subckt hw2_part2_1  VSS OUT5 VDD OUT3 OUT OUT2 IN OUT4
* 
* OUT4	OUT4
* IN	IN
* OUT2	OUT2
* OUT	OUT
* OUT3	OUT3
* VDD	VDD
* OUT5	OUT5
* VSS	VSS
MM9 N_OUT4_MM9_d N_OUT3_MM9_g N_VSS_MM9_s N_VSS_MM8_b N_18 L=1.8e-07 W=5.5e-06
+ AD=2.695e-12 AS=2.695e-12 PD=6.48e-06 PS=6.48e-06
MM11 N_OUT5_MM11_d N_OUT4_MM11_g N_VSS_MM11_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=2.695e-12 PD=5.1e-07 PS=6.48e-06
MM11@9 N_OUT5_MM11@9_d N_OUT4_MM11@9_g N_VSS_MM11@9_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@8 N_OUT5_MM11@8_d N_OUT4_MM11@8_g N_VSS_MM11@8_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@7 N_OUT5_MM11@7_d N_OUT4_MM11@7_g N_VSS_MM11@7_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@6 N_OUT5_MM11@6_d N_OUT4_MM11@6_g N_VSS_MM11@6_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@5 N_OUT5_MM11@5_d N_OUT4_MM11@5_g N_VSS_MM11@5_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@4 N_OUT5_MM11@4_d N_OUT4_MM11@4_g N_VSS_MM11@4_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@3 N_OUT5_MM11@3_d N_OUT4_MM11@3_g N_VSS_MM11@3_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=1.4025e-12 AS=1.4025e-12 PD=5.1e-07 PS=5.1e-07
MM11@2 N_OUT5_MM11@2_d N_OUT4_MM11@2_g N_VSS_MM11@2_s N_VSS_MM8_b N_18 L=1.8e-07
+ W=5.5e-06 AD=2.695e-12 AS=1.4025e-12 PD=6.48e-06 PS=5.1e-07
MM8 N_OUT3_MM8_d N_OUT2_MM8_g N_VSS_MM8_s N_VSS_MM8_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM4 N_OUT2_MM4_d N_OUT_MM4_g N_VSS_MM4_s N_VSS_MM8_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM10 N_OUT_MM10_d N_IN_MM10_g N_VSS_MM10_s N_VSS_MM8_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM7 N_OUT5_MM7_d N_OUT4_MM7_g N_VDD_MM7_s N_VDD_MM3_b P_18 L=1.8e-07 W=5e-06
+ AD=2.45e-12 AS=1.275e-12 PD=5.98e-06 PS=5.1e-07
MM7@9 N_OUT5_MM7@9_d N_OUT4_MM7@9_g N_VDD_MM7@9_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@8 N_OUT5_MM7@8_d N_OUT4_MM7@8_g N_VDD_MM7@8_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@7 N_OUT5_MM7@7_d N_OUT4_MM7@7_g N_VDD_MM7@7_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@6 N_OUT5_MM7@6_d N_OUT4_MM7@6_g N_VDD_MM7@6_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@5 N_OUT5_MM7@5_d N_OUT4_MM7@5_g N_VDD_MM7@5_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@4 N_OUT5_MM7@4_d N_OUT4_MM7@4_g N_VDD_MM7@4_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@3 N_OUT5_MM7@3_d N_OUT4_MM7@3_g N_VDD_MM7@3_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=1.275e-12 PD=5.1e-07 PS=5.1e-07
MM7@2 N_OUT5_MM7@2_d N_OUT4_MM7@2_g N_VDD_MM7@2_s N_VDD_MM3_b P_18 L=1.8e-07
+ W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
MM5 N_OUT4_MM5_d N_OUT3_MM5_g N_VDD_MM5_s N_VDD_MM3_b P_18 L=1.8e-07 W=5e-06
+ AD=2.45e-12 AS=2.45e-12 PD=5.98e-06 PS=5.98e-06
MM3 N_OUT3_MM3_d N_OUT2_MM3_g N_VDD_MM3_s N_VDD_MM3_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM0 N_OUT2_MM0_d N_OUT_MM0_g N_VDD_MM0_s N_VDD_MM3_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM6 N_OUT_MM6_d N_IN_MM6_g N_VDD_MM6_s N_VDD_MM3_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
*
.include "hw2_part2_1_smaller.pex.spi.HW2_PART2_1_SMALLER.pxi"
*
.ends
*
*
