************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: hw2_part1_2
* View Name:     schematic
* Netlisted on:  Nov  5 11:53:00 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    hw2_part1_2
* View Name:    schematic
************************************************************************

.SUBCKT hw2_part1_2 A B C OUT VDD VSS
*.PININFO A:I B:I C:I OUT:O VDD:B VSS:B
MM5 OUT C VSS VSS N_18 W=2.0u L=180.00n m=5
MM4 net5 B VSS VSS N_18 W=2.0u L=180.00n m=5
MM3 OUT A net5 VSS N_18 W=2.0u L=180.00n m=5
MM2 OUT C net21 VDD P_18 W=2.5u L=180.00n m=6
MM1 net21 B VDD VDD P_18 W=2.5u L=180.00n m=6
MM0 net21 A VDD VDD P_18 W=2.5u L=180.00n m=12
.ENDS

