* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT ROM_CELL_RANK1
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=7 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ROM_CELL_RANK1_8X2
** N=35 EP=0 IP=44 FDC=0
.ENDS
***************************************
.SUBCKT ROM_CELL_RANK1_16X16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33
** N=161 EP=33 IP=280 FDC=256
M0 18 1 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=915 $D=0
M1 18 2 34 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=2450 $D=0
M2 18 3 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=3985 $D=0
M3 18 4 50 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=5520 $D=0
M4 18 5 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=7055 $D=0
M5 18 6 66 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=8590 $D=0
M6 18 7 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=10125 $D=0
M7 18 8 82 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=11660 $D=0
M8 18 9 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=13195 $D=0
M9 18 10 98 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=14730 $D=0
M10 18 11 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=16265 $D=0
M11 18 12 114 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=17800 $D=0
M12 18 13 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=19335 $D=0
M13 18 14 130 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=20870 $D=0
M14 18 15 17 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=22405 $D=0
M15 18 16 146 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=1720 $Y=23940 $D=0
M16 35 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=915 $D=0
M17 19 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=2450 $D=0
M18 51 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=3985 $D=0
M19 19 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=5520 $D=0
M20 67 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=7055 $D=0
M21 19 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=8590 $D=0
M22 83 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=10125 $D=0
M23 19 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=11660 $D=0
M24 99 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=13195 $D=0
M25 19 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=14730 $D=0
M26 115 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=16265 $D=0
M27 19 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=17800 $D=0
M28 131 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=19335 $D=0
M29 19 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=20870 $D=0
M30 147 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=22405 $D=0
M31 19 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=2410 $Y=23940 $D=0
M32 18 1 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=915 $D=0
M33 18 2 36 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=2450 $D=0
M34 18 3 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=3985 $D=0
M35 18 4 52 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=5520 $D=0
M36 18 5 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=7055 $D=0
M37 18 6 68 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=8590 $D=0
M38 18 7 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=10125 $D=0
M39 18 8 84 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=11660 $D=0
M40 18 9 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=13195 $D=0
M41 18 10 100 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=14730 $D=0
M42 18 11 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=16265 $D=0
M43 18 12 116 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=17800 $D=0
M44 18 13 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=19335 $D=0
M45 18 14 132 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=20870 $D=0
M46 18 15 20 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=22405 $D=0
M47 18 16 148 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=3870 $Y=23940 $D=0
M48 37 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=915 $D=0
M49 21 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=2450 $D=0
M50 53 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=3985 $D=0
M51 21 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=5520 $D=0
M52 69 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=7055 $D=0
M53 21 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=8590 $D=0
M54 85 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=10125 $D=0
M55 21 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=11660 $D=0
M56 101 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=13195 $D=0
M57 21 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=14730 $D=0
M58 117 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=16265 $D=0
M59 21 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=17800 $D=0
M60 133 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=19335 $D=0
M61 21 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=20870 $D=0
M62 149 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=22405 $D=0
M63 21 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=4560 $Y=23940 $D=0
M64 18 1 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=915 $D=0
M65 18 2 38 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=2450 $D=0
M66 18 3 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=3985 $D=0
M67 18 4 54 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=5520 $D=0
M68 18 5 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=7055 $D=0
M69 18 6 70 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=8590 $D=0
M70 18 7 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=10125 $D=0
M71 18 8 86 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=11660 $D=0
M72 18 9 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=13195 $D=0
M73 18 10 102 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=14730 $D=0
M74 18 11 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=16265 $D=0
M75 18 12 118 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=17800 $D=0
M76 18 13 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=19335 $D=0
M77 18 14 134 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=20870 $D=0
M78 18 15 22 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=22405 $D=0
M79 18 16 150 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=6020 $Y=23940 $D=0
M80 39 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=915 $D=0
M81 23 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=2450 $D=0
M82 55 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=3985 $D=0
M83 23 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=5520 $D=0
M84 71 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=7055 $D=0
M85 23 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=8590 $D=0
M86 87 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=10125 $D=0
M87 23 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=11660 $D=0
M88 103 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=13195 $D=0
M89 23 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=14730 $D=0
M90 119 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=16265 $D=0
M91 23 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=17800 $D=0
M92 135 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=19335 $D=0
M93 23 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=20870 $D=0
M94 151 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=22405 $D=0
M95 23 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=6710 $Y=23940 $D=0
M96 18 1 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=915 $D=0
M97 18 2 40 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=2450 $D=0
M98 18 3 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=3985 $D=0
M99 18 4 56 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=5520 $D=0
M100 18 5 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=7055 $D=0
M101 18 6 72 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=8590 $D=0
M102 18 7 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=10125 $D=0
M103 18 8 88 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=11660 $D=0
M104 18 9 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=13195 $D=0
M105 18 10 104 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=14730 $D=0
M106 18 11 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=16265 $D=0
M107 18 12 120 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=17800 $D=0
M108 18 13 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=19335 $D=0
M109 18 14 136 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=20870 $D=0
M110 18 15 24 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=22405 $D=0
M111 18 16 152 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=8170 $Y=23940 $D=0
M112 41 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=915 $D=0
M113 25 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=2450 $D=0
M114 57 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=3985 $D=0
M115 25 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=5520 $D=0
M116 73 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=7055 $D=0
M117 25 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=8590 $D=0
M118 89 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=10125 $D=0
M119 25 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=11660 $D=0
M120 105 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=13195 $D=0
M121 25 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=14730 $D=0
M122 121 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=16265 $D=0
M123 25 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=17800 $D=0
M124 137 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=19335 $D=0
M125 25 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=20870 $D=0
M126 153 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=22405 $D=0
M127 25 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=8860 $Y=23940 $D=0
M128 18 1 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=915 $D=0
M129 18 2 42 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=2450 $D=0
M130 18 3 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=3985 $D=0
M131 18 4 58 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=5520 $D=0
M132 18 5 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=7055 $D=0
M133 18 6 74 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=8590 $D=0
M134 18 7 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=10125 $D=0
M135 18 8 90 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=11660 $D=0
M136 18 9 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=13195 $D=0
M137 18 10 106 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=14730 $D=0
M138 18 11 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=16265 $D=0
M139 18 12 122 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=17800 $D=0
M140 18 13 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=19335 $D=0
M141 18 14 138 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=20870 $D=0
M142 18 15 26 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=22405 $D=0
M143 18 16 154 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=10320 $Y=23940 $D=0
M144 43 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=915 $D=0
M145 27 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=2450 $D=0
M146 59 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=3985 $D=0
M147 27 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=5520 $D=0
M148 75 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=7055 $D=0
M149 27 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=8590 $D=0
M150 91 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=10125 $D=0
M151 27 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=11660 $D=0
M152 107 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=13195 $D=0
M153 27 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=14730 $D=0
M154 123 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=16265 $D=0
M155 27 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=17800 $D=0
M156 139 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=19335 $D=0
M157 27 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=20870 $D=0
M158 155 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=22405 $D=0
M159 27 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=11010 $Y=23940 $D=0
M160 18 1 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=915 $D=0
M161 18 2 44 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=2450 $D=0
M162 18 3 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=3985 $D=0
M163 18 4 60 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=5520 $D=0
M164 18 5 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=7055 $D=0
M165 18 6 76 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=8590 $D=0
M166 18 7 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=10125 $D=0
M167 18 8 92 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=11660 $D=0
M168 18 9 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=13195 $D=0
M169 18 10 108 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=14730 $D=0
M170 18 11 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=16265 $D=0
M171 18 12 124 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=17800 $D=0
M172 18 13 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=19335 $D=0
M173 18 14 140 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=20870 $D=0
M174 18 15 28 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=22405 $D=0
M175 18 16 156 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=12470 $Y=23940 $D=0
M176 45 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=915 $D=0
M177 29 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=2450 $D=0
M178 61 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=3985 $D=0
M179 29 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=5520 $D=0
M180 77 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=7055 $D=0
M181 29 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=8590 $D=0
M182 93 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=10125 $D=0
M183 29 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=11660 $D=0
M184 109 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=13195 $D=0
M185 29 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=14730 $D=0
M186 125 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=16265 $D=0
M187 29 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=17800 $D=0
M188 141 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=19335 $D=0
M189 29 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=20870 $D=0
M190 157 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=22405 $D=0
M191 29 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=13160 $Y=23940 $D=0
M192 18 1 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=915 $D=0
M193 18 2 46 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=2450 $D=0
M194 18 3 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=3985 $D=0
M195 18 4 62 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=5520 $D=0
M196 18 5 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=7055 $D=0
M197 18 6 78 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=8590 $D=0
M198 18 7 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=10125 $D=0
M199 18 8 94 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=11660 $D=0
M200 18 9 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=13195 $D=0
M201 18 10 110 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=14730 $D=0
M202 18 11 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=16265 $D=0
M203 18 12 126 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=17800 $D=0
M204 18 13 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=19335 $D=0
M205 18 14 142 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=20870 $D=0
M206 18 15 30 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=22405 $D=0
M207 18 16 158 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=14620 $Y=23940 $D=0
M208 47 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=915 $D=0
M209 31 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=2450 $D=0
M210 63 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=3985 $D=0
M211 31 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=5520 $D=0
M212 79 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=7055 $D=0
M213 31 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=8590 $D=0
M214 95 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=10125 $D=0
M215 31 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=11660 $D=0
M216 111 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=13195 $D=0
M217 31 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=14730 $D=0
M218 127 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=16265 $D=0
M219 31 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=17800 $D=0
M220 143 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=19335 $D=0
M221 31 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=20870 $D=0
M222 159 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=22405 $D=0
M223 31 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=15310 $Y=23940 $D=0
M224 18 1 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=915 $D=0
M225 18 2 48 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=2450 $D=0
M226 18 3 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=3985 $D=0
M227 18 4 64 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=5520 $D=0
M228 18 5 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=7055 $D=0
M229 18 6 80 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=8590 $D=0
M230 18 7 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=10125 $D=0
M231 18 8 96 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=11660 $D=0
M232 18 9 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=13195 $D=0
M233 18 10 112 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=14730 $D=0
M234 18 11 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=16265 $D=0
M235 18 12 128 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=17800 $D=0
M236 18 13 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=19335 $D=0
M237 18 14 144 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=20870 $D=0
M238 18 15 32 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=22405 $D=0
M239 18 16 160 18 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=16770 $Y=23940 $D=0
M240 49 1 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=915 $D=0
M241 33 2 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=2450 $D=0
M242 65 3 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=3985 $D=0
M243 33 4 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=5520 $D=0
M244 81 5 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=7055 $D=0
M245 33 6 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=8590 $D=0
M246 97 7 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=10125 $D=0
M247 33 8 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=11660 $D=0
M248 113 9 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=13195 $D=0
M249 33 10 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=14730 $D=0
M250 129 11 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=16265 $D=0
M251 33 12 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=17800 $D=0
M252 145 13 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=19335 $D=0
M253 33 14 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=20870 $D=0
M254 161 15 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=22405 $D=0
M255 33 16 18 18 N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=17460 $Y=23940 $D=0
.ENDS
***************************************
.SUBCKT ROM_CELL_RANK1_16X64 BL<0> VSS BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15> WL<63> WL<47> WL<31>
+ WL<15> WL<62> WL<46> WL<30> WL<14> WL<61> WL<45> WL<29> WL<13> WL<60> WL<44> WL<28> WL<12> WL<59> WL<43> WL<27> WL<11> WL<58> WL<42> WL<26>
+ WL<10> WL<57> WL<41> WL<25> WL<9> WL<56> WL<40> WL<24> WL<8> WL<55> WL<39> WL<23> WL<7> WL<54> WL<38> WL<22> WL<6> WL<53> WL<37> WL<21>
+ WL<5> WL<52> WL<36> WL<20> WL<4> WL<51> WL<35> WL<19> WL<3> WL<50> WL<34> WL<18> WL<2> WL<49> WL<33> WL<17> WL<1> WL<48> WL<32> WL<16>
+ WL<0>
** N=81 EP=81 IP=132 FDC=1024
X0 WL<63> WL<62> WL<61> WL<60> WL<59> WL<58> WL<57> WL<56> WL<55> WL<54> WL<53> WL<52> WL<51> WL<50> WL<49> WL<48> BL<0> VSS BL<1> BL<2>
+ BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15>
+ ROM_CELL_RANK1_16X16 $T=0 0 0 0 $X=0 $Y=0
X1 WL<47> WL<46> WL<45> WL<44> WL<43> WL<42> WL<41> WL<40> WL<39> WL<38> WL<37> WL<36> WL<35> WL<34> WL<33> WL<32> BL<0> VSS BL<1> BL<2>
+ BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15>
+ ROM_CELL_RANK1_16X16 $T=0 24980 0 0 $X=0 $Y=24980
X2 WL<31> WL<30> WL<29> WL<28> WL<27> WL<26> WL<25> WL<24> WL<23> WL<22> WL<21> WL<20> WL<19> WL<18> WL<17> WL<16> BL<0> VSS BL<1> BL<2>
+ BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15>
+ ROM_CELL_RANK1_16X16 $T=0 49960 0 0 $X=0 $Y=49960
X3 WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0> BL<0> VSS BL<1> BL<2>
+ BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15>
+ ROM_CELL_RANK1_16X16 $T=0 74940 0 0 $X=0 $Y=74940
.ENDS
***************************************
