* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT final_precharge WL<63> WL<62> WL<61> WL<60> WL<59> WL<58> WL<57> WL<56> WL<55> WL<54> WL<53> WL<52> WL<51> WL<50> WL<49> WL<48> WL<47> WL<46> WL<45> WL<44>
+ WL<43> WL<42> WL<41> WL<40> WL<39> WL<38> WL<37> WL<36> WL<35> WL<34> WL<33> WL<32> WL<31> WL<30> WL<29> WL<28> WL<27> WL<26> WL<25> WL<24>
+ WL<23> WL<22> WL<21> WL<20> WL<19> WL<18> WL<17> WL<16> WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> WL<9> WL<8> WL<7> WL<6> WL<5> WL<4>
+ WL<3> WL<2> WL<1> WL<0> BL<0> VSS BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14>
+ pre_b BL<15> VDD
** N=595 EP=83 IP=0 FDC=1040
M0 VSS WL<63> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-37140 $D=0
M1 VSS WL<62> 83 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-35605 $D=0
M2 VSS WL<61> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-34070 $D=0
M3 VSS WL<60> 84 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-32535 $D=0
M4 VSS WL<59> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-31000 $D=0
M5 VSS WL<58> 85 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-29465 $D=0
M6 VSS WL<57> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-27930 $D=0
M7 VSS WL<56> 86 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-26395 $D=0
M8 VSS WL<55> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-24860 $D=0
M9 VSS WL<54> 87 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-23325 $D=0
M10 VSS WL<53> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-21790 $D=0
M11 VSS WL<52> 88 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-20255 $D=0
M12 VSS WL<51> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-18720 $D=0
M13 VSS WL<50> 89 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-17185 $D=0
M14 VSS WL<49> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-15650 $D=0
M15 VSS WL<48> 90 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-14115 $D=0
M16 VSS WL<47> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-12160 $D=0
M17 VSS WL<46> 91 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-10625 $D=0
M18 VSS WL<45> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-9090 $D=0
M19 VSS WL<44> 92 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-7555 $D=0
M20 VSS WL<43> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-6020 $D=0
M21 VSS WL<42> 93 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-4485 $D=0
M22 VSS WL<41> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-2950 $D=0
M23 VSS WL<40> 94 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=-1415 $D=0
M24 VSS WL<39> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=120 $D=0
M25 VSS WL<38> 95 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=1655 $D=0
M26 VSS WL<37> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=3190 $D=0
M27 VSS WL<36> 96 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=4725 $D=0
M28 VSS WL<35> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=6260 $D=0
M29 VSS WL<34> 97 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=7795 $D=0
M30 VSS WL<33> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=9330 $D=0
M31 VSS WL<32> 98 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=10865 $D=0
M32 VSS WL<31> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=12820 $D=0
M33 VSS WL<30> 99 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=14355 $D=0
M34 VSS WL<29> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=15890 $D=0
M35 VSS WL<28> 100 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=17425 $D=0
M36 VSS WL<27> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=18960 $D=0
M37 VSS WL<26> 101 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=20495 $D=0
M38 VSS WL<25> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=22030 $D=0
M39 VSS WL<24> 102 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=23565 $D=0
M40 VSS WL<23> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=25100 $D=0
M41 VSS WL<22> 103 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=26635 $D=0
M42 VSS WL<21> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=28170 $D=0
M43 VSS WL<20> 104 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=29705 $D=0
M44 VSS WL<19> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=31240 $D=0
M45 VSS WL<18> 105 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=32775 $D=0
M46 VSS WL<17> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=34310 $D=0
M47 VSS WL<16> 106 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=35845 $D=0
M48 VSS WL<15> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=37800 $D=0
M49 VSS WL<14> 107 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=39335 $D=0
M50 VSS WL<13> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=40870 $D=0
M51 VSS WL<12> 108 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=42405 $D=0
M52 VSS WL<11> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=43940 $D=0
M53 VSS WL<10> 109 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=45475 $D=0
M54 VSS WL<9> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=47010 $D=0
M55 VSS WL<8> 110 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=48545 $D=0
M56 VSS WL<7> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=50080 $D=0
M57 VSS WL<6> 111 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=51615 $D=0
M58 VSS WL<5> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=53150 $D=0
M59 VSS WL<4> 112 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=54685 $D=0
M60 VSS WL<3> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=56220 $D=0
M61 VSS WL<2> 113 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=57755 $D=0
M62 VSS WL<1> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=59290 $D=0
M63 VSS WL<0> 114 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=24085 $Y=60825 $D=0
M64 115 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-37140 $D=0
M65 BL<1> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-35605 $D=0
M66 116 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-34070 $D=0
M67 BL<1> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-32535 $D=0
M68 117 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-31000 $D=0
M69 BL<1> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-29465 $D=0
M70 118 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-27930 $D=0
M71 BL<1> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-26395 $D=0
M72 119 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-24860 $D=0
M73 BL<1> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-23325 $D=0
M74 120 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-21790 $D=0
M75 BL<1> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-20255 $D=0
M76 121 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-18720 $D=0
M77 BL<1> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-17185 $D=0
M78 122 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-15650 $D=0
M79 BL<1> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-14115 $D=0
M80 123 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-12160 $D=0
M81 BL<1> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-10625 $D=0
M82 124 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-9090 $D=0
M83 BL<1> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-7555 $D=0
M84 125 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-6020 $D=0
M85 BL<1> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-4485 $D=0
M86 126 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-2950 $D=0
M87 BL<1> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=-1415 $D=0
M88 127 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=120 $D=0
M89 BL<1> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=1655 $D=0
M90 128 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=3190 $D=0
M91 BL<1> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=4725 $D=0
M92 129 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=6260 $D=0
M93 BL<1> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=7795 $D=0
M94 130 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=9330 $D=0
M95 BL<1> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=10865 $D=0
M96 131 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=12820 $D=0
M97 BL<1> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=14355 $D=0
M98 132 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=15890 $D=0
M99 BL<1> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=17425 $D=0
M100 133 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=18960 $D=0
M101 BL<1> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=20495 $D=0
M102 134 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=22030 $D=0
M103 BL<1> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=23565 $D=0
M104 135 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=25100 $D=0
M105 BL<1> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=26635 $D=0
M106 136 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=28170 $D=0
M107 BL<1> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=29705 $D=0
M108 137 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=31240 $D=0
M109 BL<1> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=32775 $D=0
M110 138 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=34310 $D=0
M111 BL<1> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=35845 $D=0
M112 139 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=37800 $D=0
M113 BL<1> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=39335 $D=0
M114 140 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=40870 $D=0
M115 BL<1> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=42405 $D=0
M116 141 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=43940 $D=0
M117 BL<1> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=45475 $D=0
M118 142 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=47010 $D=0
M119 BL<1> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=48545 $D=0
M120 143 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=50080 $D=0
M121 BL<1> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=51615 $D=0
M122 144 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=53150 $D=0
M123 BL<1> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=54685 $D=0
M124 145 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=56220 $D=0
M125 BL<1> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=57755 $D=0
M126 146 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=59290 $D=0
M127 BL<1> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=24775 $Y=60825 $D=0
M128 VSS WL<63> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-37140 $D=0
M129 VSS WL<62> 147 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-35605 $D=0
M130 VSS WL<61> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-34070 $D=0
M131 VSS WL<60> 148 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-32535 $D=0
M132 VSS WL<59> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-31000 $D=0
M133 VSS WL<58> 149 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-29465 $D=0
M134 VSS WL<57> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-27930 $D=0
M135 VSS WL<56> 150 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-26395 $D=0
M136 VSS WL<55> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-24860 $D=0
M137 VSS WL<54> 151 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-23325 $D=0
M138 VSS WL<53> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-21790 $D=0
M139 VSS WL<52> 152 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-20255 $D=0
M140 VSS WL<51> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-18720 $D=0
M141 VSS WL<50> 153 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-17185 $D=0
M142 VSS WL<49> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-15650 $D=0
M143 VSS WL<48> 154 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-14115 $D=0
M144 VSS WL<47> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-12160 $D=0
M145 VSS WL<46> 155 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-10625 $D=0
M146 VSS WL<45> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-9090 $D=0
M147 VSS WL<44> 156 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-7555 $D=0
M148 VSS WL<43> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-6020 $D=0
M149 VSS WL<42> 157 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-4485 $D=0
M150 VSS WL<41> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-2950 $D=0
M151 VSS WL<40> 158 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=-1415 $D=0
M152 VSS WL<39> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=120 $D=0
M153 VSS WL<38> 159 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=1655 $D=0
M154 VSS WL<37> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=3190 $D=0
M155 VSS WL<36> 160 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=4725 $D=0
M156 VSS WL<35> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=6260 $D=0
M157 VSS WL<34> 161 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=7795 $D=0
M158 VSS WL<33> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=9330 $D=0
M159 VSS WL<32> 162 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=10865 $D=0
M160 VSS WL<31> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=12820 $D=0
M161 VSS WL<30> 163 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=14355 $D=0
M162 VSS WL<29> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=15890 $D=0
M163 VSS WL<28> 164 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=17425 $D=0
M164 VSS WL<27> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=18960 $D=0
M165 VSS WL<26> 165 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=20495 $D=0
M166 VSS WL<25> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=22030 $D=0
M167 VSS WL<24> 166 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=23565 $D=0
M168 VSS WL<23> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=25100 $D=0
M169 VSS WL<22> 167 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=26635 $D=0
M170 VSS WL<21> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=28170 $D=0
M171 VSS WL<20> 168 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=29705 $D=0
M172 VSS WL<19> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=31240 $D=0
M173 VSS WL<18> 169 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=32775 $D=0
M174 VSS WL<17> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=34310 $D=0
M175 VSS WL<16> 170 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=35845 $D=0
M176 VSS WL<15> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=37800 $D=0
M177 VSS WL<14> 171 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=39335 $D=0
M178 VSS WL<13> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=40870 $D=0
M179 VSS WL<12> 172 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=42405 $D=0
M180 VSS WL<11> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=43940 $D=0
M181 VSS WL<10> 173 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=45475 $D=0
M182 VSS WL<9> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=47010 $D=0
M183 VSS WL<8> 174 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=48545 $D=0
M184 VSS WL<7> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=50080 $D=0
M185 VSS WL<6> 175 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=51615 $D=0
M186 VSS WL<5> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=53150 $D=0
M187 VSS WL<4> 176 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=54685 $D=0
M188 VSS WL<3> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=56220 $D=0
M189 VSS WL<2> 177 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=57755 $D=0
M190 VSS WL<1> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=59290 $D=0
M191 VSS WL<0> 178 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=26235 $Y=60825 $D=0
M192 179 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-37140 $D=0
M193 BL<3> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-35605 $D=0
M194 180 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-34070 $D=0
M195 BL<3> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-32535 $D=0
M196 181 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-31000 $D=0
M197 BL<3> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-29465 $D=0
M198 182 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-27930 $D=0
M199 BL<3> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-26395 $D=0
M200 183 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-24860 $D=0
M201 BL<3> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-23325 $D=0
M202 184 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-21790 $D=0
M203 BL<3> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-20255 $D=0
M204 185 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-18720 $D=0
M205 BL<3> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-17185 $D=0
M206 186 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-15650 $D=0
M207 BL<3> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-14115 $D=0
M208 187 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-12160 $D=0
M209 BL<3> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-10625 $D=0
M210 188 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-9090 $D=0
M211 BL<3> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-7555 $D=0
M212 189 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-6020 $D=0
M213 BL<3> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-4485 $D=0
M214 190 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-2950 $D=0
M215 BL<3> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=-1415 $D=0
M216 191 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=120 $D=0
M217 BL<3> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=1655 $D=0
M218 192 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=3190 $D=0
M219 BL<3> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=4725 $D=0
M220 193 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=6260 $D=0
M221 BL<3> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=7795 $D=0
M222 194 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=9330 $D=0
M223 BL<3> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=10865 $D=0
M224 195 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=12820 $D=0
M225 BL<3> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=14355 $D=0
M226 196 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=15890 $D=0
M227 BL<3> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=17425 $D=0
M228 197 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=18960 $D=0
M229 BL<3> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=20495 $D=0
M230 198 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=22030 $D=0
M231 BL<3> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=23565 $D=0
M232 199 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=25100 $D=0
M233 BL<3> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=26635 $D=0
M234 200 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=28170 $D=0
M235 BL<3> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=29705 $D=0
M236 201 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=31240 $D=0
M237 BL<3> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=32775 $D=0
M238 202 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=34310 $D=0
M239 BL<3> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=35845 $D=0
M240 203 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=37800 $D=0
M241 BL<3> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=39335 $D=0
M242 204 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=40870 $D=0
M243 BL<3> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=42405 $D=0
M244 205 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=43940 $D=0
M245 BL<3> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=45475 $D=0
M246 206 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=47010 $D=0
M247 BL<3> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=48545 $D=0
M248 207 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=50080 $D=0
M249 BL<3> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=51615 $D=0
M250 208 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=53150 $D=0
M251 BL<3> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=54685 $D=0
M252 209 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=56220 $D=0
M253 BL<3> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=57755 $D=0
M254 210 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=59290 $D=0
M255 BL<3> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=26925 $Y=60825 $D=0
M256 VSS WL<63> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-37140 $D=0
M257 VSS WL<62> 211 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-35605 $D=0
M258 VSS WL<61> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-34070 $D=0
M259 VSS WL<60> 212 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-32535 $D=0
M260 VSS WL<59> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-31000 $D=0
M261 VSS WL<58> 213 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-29465 $D=0
M262 VSS WL<57> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-27930 $D=0
M263 VSS WL<56> 214 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-26395 $D=0
M264 VSS WL<55> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-24860 $D=0
M265 VSS WL<54> 215 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-23325 $D=0
M266 VSS WL<53> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-21790 $D=0
M267 VSS WL<52> 216 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-20255 $D=0
M268 VSS WL<51> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-18720 $D=0
M269 VSS WL<50> 217 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-17185 $D=0
M270 VSS WL<49> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-15650 $D=0
M271 VSS WL<48> 218 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-14115 $D=0
M272 VSS WL<47> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-12160 $D=0
M273 VSS WL<46> 219 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-10625 $D=0
M274 VSS WL<45> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-9090 $D=0
M275 VSS WL<44> 220 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-7555 $D=0
M276 VSS WL<43> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-6020 $D=0
M277 VSS WL<42> 221 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-4485 $D=0
M278 VSS WL<41> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-2950 $D=0
M279 VSS WL<40> 222 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=-1415 $D=0
M280 VSS WL<39> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=120 $D=0
M281 VSS WL<38> 223 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=1655 $D=0
M282 VSS WL<37> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=3190 $D=0
M283 VSS WL<36> 224 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=4725 $D=0
M284 VSS WL<35> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=6260 $D=0
M285 VSS WL<34> 225 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=7795 $D=0
M286 VSS WL<33> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=9330 $D=0
M287 VSS WL<32> 226 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=10865 $D=0
M288 VSS WL<31> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=12820 $D=0
M289 VSS WL<30> 227 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=14355 $D=0
M290 VSS WL<29> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=15890 $D=0
M291 VSS WL<28> 228 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=17425 $D=0
M292 VSS WL<27> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=18960 $D=0
M293 VSS WL<26> 229 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=20495 $D=0
M294 VSS WL<25> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=22030 $D=0
M295 VSS WL<24> 230 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=23565 $D=0
M296 VSS WL<23> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=25100 $D=0
M297 VSS WL<22> 231 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=26635 $D=0
M298 VSS WL<21> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=28170 $D=0
M299 VSS WL<20> 232 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=29705 $D=0
M300 VSS WL<19> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=31240 $D=0
M301 VSS WL<18> 233 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=32775 $D=0
M302 VSS WL<17> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=34310 $D=0
M303 VSS WL<16> 234 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=35845 $D=0
M304 VSS WL<15> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=37800 $D=0
M305 VSS WL<14> 235 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=39335 $D=0
M306 VSS WL<13> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=40870 $D=0
M307 VSS WL<12> 236 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=42405 $D=0
M308 VSS WL<11> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=43940 $D=0
M309 VSS WL<10> 237 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=45475 $D=0
M310 VSS WL<9> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=47010 $D=0
M311 VSS WL<8> 238 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=48545 $D=0
M312 VSS WL<7> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=50080 $D=0
M313 VSS WL<6> 239 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=51615 $D=0
M314 VSS WL<5> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=53150 $D=0
M315 VSS WL<4> 240 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=54685 $D=0
M316 VSS WL<3> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=56220 $D=0
M317 VSS WL<2> 241 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=57755 $D=0
M318 VSS WL<1> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=59290 $D=0
M319 VSS WL<0> 242 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=28385 $Y=60825 $D=0
M320 243 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-37140 $D=0
M321 BL<5> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-35605 $D=0
M322 244 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-34070 $D=0
M323 BL<5> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-32535 $D=0
M324 245 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-31000 $D=0
M325 BL<5> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-29465 $D=0
M326 246 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-27930 $D=0
M327 BL<5> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-26395 $D=0
M328 247 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-24860 $D=0
M329 BL<5> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-23325 $D=0
M330 248 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-21790 $D=0
M331 BL<5> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-20255 $D=0
M332 249 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-18720 $D=0
M333 BL<5> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-17185 $D=0
M334 250 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-15650 $D=0
M335 BL<5> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-14115 $D=0
M336 251 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-12160 $D=0
M337 BL<5> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-10625 $D=0
M338 252 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-9090 $D=0
M339 BL<5> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-7555 $D=0
M340 253 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-6020 $D=0
M341 BL<5> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-4485 $D=0
M342 254 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-2950 $D=0
M343 BL<5> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=-1415 $D=0
M344 255 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=120 $D=0
M345 BL<5> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=1655 $D=0
M346 256 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=3190 $D=0
M347 BL<5> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=4725 $D=0
M348 257 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=6260 $D=0
M349 BL<5> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=7795 $D=0
M350 258 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=9330 $D=0
M351 BL<5> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=10865 $D=0
M352 259 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=12820 $D=0
M353 BL<5> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=14355 $D=0
M354 260 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=15890 $D=0
M355 BL<5> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=17425 $D=0
M356 261 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=18960 $D=0
M357 BL<5> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=20495 $D=0
M358 262 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=22030 $D=0
M359 BL<5> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=23565 $D=0
M360 263 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=25100 $D=0
M361 BL<5> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=26635 $D=0
M362 264 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=28170 $D=0
M363 BL<5> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=29705 $D=0
M364 265 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=31240 $D=0
M365 BL<5> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=32775 $D=0
M366 266 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=34310 $D=0
M367 BL<5> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=35845 $D=0
M368 267 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=37800 $D=0
M369 BL<5> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=39335 $D=0
M370 268 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=40870 $D=0
M371 BL<5> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=42405 $D=0
M372 269 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=43940 $D=0
M373 BL<5> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=45475 $D=0
M374 270 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=47010 $D=0
M375 BL<5> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=48545 $D=0
M376 271 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=50080 $D=0
M377 BL<5> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=51615 $D=0
M378 272 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=53150 $D=0
M379 BL<5> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=54685 $D=0
M380 273 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=56220 $D=0
M381 BL<5> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=57755 $D=0
M382 274 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=59290 $D=0
M383 BL<5> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=29075 $Y=60825 $D=0
M384 VSS WL<63> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-37140 $D=0
M385 VSS WL<62> 275 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-35605 $D=0
M386 VSS WL<61> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-34070 $D=0
M387 VSS WL<60> 276 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-32535 $D=0
M388 VSS WL<59> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-31000 $D=0
M389 VSS WL<58> 277 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-29465 $D=0
M390 VSS WL<57> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-27930 $D=0
M391 VSS WL<56> 278 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-26395 $D=0
M392 VSS WL<55> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-24860 $D=0
M393 VSS WL<54> 279 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-23325 $D=0
M394 VSS WL<53> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-21790 $D=0
M395 VSS WL<52> 280 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-20255 $D=0
M396 VSS WL<51> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-18720 $D=0
M397 VSS WL<50> 281 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-17185 $D=0
M398 VSS WL<49> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-15650 $D=0
M399 VSS WL<48> 282 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-14115 $D=0
M400 VSS WL<47> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-12160 $D=0
M401 VSS WL<46> 283 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-10625 $D=0
M402 VSS WL<45> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-9090 $D=0
M403 VSS WL<44> 284 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-7555 $D=0
M404 VSS WL<43> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-6020 $D=0
M405 VSS WL<42> 285 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-4485 $D=0
M406 VSS WL<41> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-2950 $D=0
M407 VSS WL<40> 286 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=-1415 $D=0
M408 VSS WL<39> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=120 $D=0
M409 VSS WL<38> 287 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=1655 $D=0
M410 VSS WL<37> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=3190 $D=0
M411 VSS WL<36> 288 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=4725 $D=0
M412 VSS WL<35> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=6260 $D=0
M413 VSS WL<34> 289 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=7795 $D=0
M414 VSS WL<33> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=9330 $D=0
M415 VSS WL<32> 290 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=10865 $D=0
M416 VSS WL<31> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=12820 $D=0
M417 VSS WL<30> 291 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=14355 $D=0
M418 VSS WL<29> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=15890 $D=0
M419 VSS WL<28> 292 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=17425 $D=0
M420 VSS WL<27> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=18960 $D=0
M421 VSS WL<26> 293 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=20495 $D=0
M422 VSS WL<25> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=22030 $D=0
M423 VSS WL<24> 294 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=23565 $D=0
M424 VSS WL<23> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=25100 $D=0
M425 VSS WL<22> 295 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=26635 $D=0
M426 VSS WL<21> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=28170 $D=0
M427 VSS WL<20> 296 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=29705 $D=0
M428 VSS WL<19> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=31240 $D=0
M429 VSS WL<18> 297 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=32775 $D=0
M430 VSS WL<17> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=34310 $D=0
M431 VSS WL<16> 298 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=35845 $D=0
M432 VSS WL<15> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=37800 $D=0
M433 VSS WL<14> 299 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=39335 $D=0
M434 VSS WL<13> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=40870 $D=0
M435 VSS WL<12> 300 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=42405 $D=0
M436 VSS WL<11> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=43940 $D=0
M437 VSS WL<10> 301 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=45475 $D=0
M438 VSS WL<9> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=47010 $D=0
M439 VSS WL<8> 302 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=48545 $D=0
M440 VSS WL<7> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=50080 $D=0
M441 VSS WL<6> 303 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=51615 $D=0
M442 VSS WL<5> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=53150 $D=0
M443 VSS WL<4> 304 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=54685 $D=0
M444 VSS WL<3> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=56220 $D=0
M445 VSS WL<2> 305 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=57755 $D=0
M446 VSS WL<1> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=59290 $D=0
M447 VSS WL<0> 306 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=30535 $Y=60825 $D=0
M448 307 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-37140 $D=0
M449 BL<7> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-35605 $D=0
M450 308 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-34070 $D=0
M451 BL<7> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-32535 $D=0
M452 309 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-31000 $D=0
M453 BL<7> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-29465 $D=0
M454 310 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-27930 $D=0
M455 BL<7> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-26395 $D=0
M456 311 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-24860 $D=0
M457 BL<7> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-23325 $D=0
M458 312 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-21790 $D=0
M459 BL<7> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-20255 $D=0
M460 313 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-18720 $D=0
M461 BL<7> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-17185 $D=0
M462 314 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-15650 $D=0
M463 BL<7> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-14115 $D=0
M464 315 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-12160 $D=0
M465 BL<7> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-10625 $D=0
M466 316 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-9090 $D=0
M467 BL<7> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-7555 $D=0
M468 317 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-6020 $D=0
M469 BL<7> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-4485 $D=0
M470 318 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-2950 $D=0
M471 BL<7> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=-1415 $D=0
M472 319 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=120 $D=0
M473 BL<7> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=1655 $D=0
M474 320 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=3190 $D=0
M475 BL<7> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=4725 $D=0
M476 321 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=6260 $D=0
M477 BL<7> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=7795 $D=0
M478 322 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=9330 $D=0
M479 BL<7> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=10865 $D=0
M480 323 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=12820 $D=0
M481 BL<7> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=14355 $D=0
M482 324 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=15890 $D=0
M483 BL<7> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=17425 $D=0
M484 325 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=18960 $D=0
M485 BL<7> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=20495 $D=0
M486 326 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=22030 $D=0
M487 BL<7> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=23565 $D=0
M488 327 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=25100 $D=0
M489 BL<7> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=26635 $D=0
M490 328 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=28170 $D=0
M491 BL<7> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=29705 $D=0
M492 329 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=31240 $D=0
M493 BL<7> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=32775 $D=0
M494 330 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=34310 $D=0
M495 BL<7> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=35845 $D=0
M496 331 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=37800 $D=0
M497 BL<7> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=39335 $D=0
M498 332 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=40870 $D=0
M499 BL<7> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=42405 $D=0
M500 333 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=43940 $D=0
M501 BL<7> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=45475 $D=0
M502 334 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=47010 $D=0
M503 BL<7> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=48545 $D=0
M504 335 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=50080 $D=0
M505 BL<7> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=51615 $D=0
M506 336 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=53150 $D=0
M507 BL<7> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=54685 $D=0
M508 337 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=56220 $D=0
M509 BL<7> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=57755 $D=0
M510 338 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=59290 $D=0
M511 BL<7> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=31225 $Y=60825 $D=0
M512 VSS WL<63> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-37140 $D=0
M513 VSS WL<62> 339 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-35605 $D=0
M514 VSS WL<61> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-34070 $D=0
M515 VSS WL<60> 340 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-32535 $D=0
M516 VSS WL<59> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-31000 $D=0
M517 VSS WL<58> 341 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-29465 $D=0
M518 VSS WL<57> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-27930 $D=0
M519 VSS WL<56> 342 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-26395 $D=0
M520 VSS WL<55> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-24860 $D=0
M521 VSS WL<54> 343 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-23325 $D=0
M522 VSS WL<53> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-21790 $D=0
M523 VSS WL<52> 344 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-20255 $D=0
M524 VSS WL<51> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-18720 $D=0
M525 VSS WL<50> 345 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-17185 $D=0
M526 VSS WL<49> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-15650 $D=0
M527 VSS WL<48> 346 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-14115 $D=0
M528 VSS WL<47> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-12160 $D=0
M529 VSS WL<46> 347 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-10625 $D=0
M530 VSS WL<45> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-9090 $D=0
M531 VSS WL<44> 348 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-7555 $D=0
M532 VSS WL<43> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-6020 $D=0
M533 VSS WL<42> 349 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-4485 $D=0
M534 VSS WL<41> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-2950 $D=0
M535 VSS WL<40> 350 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=-1415 $D=0
M536 VSS WL<39> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=120 $D=0
M537 VSS WL<38> 351 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=1655 $D=0
M538 VSS WL<37> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=3190 $D=0
M539 VSS WL<36> 352 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=4725 $D=0
M540 VSS WL<35> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=6260 $D=0
M541 VSS WL<34> 353 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=7795 $D=0
M542 VSS WL<33> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=9330 $D=0
M543 VSS WL<32> 354 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=10865 $D=0
M544 VSS WL<31> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=12820 $D=0
M545 VSS WL<30> 355 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=14355 $D=0
M546 VSS WL<29> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=15890 $D=0
M547 VSS WL<28> 356 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=17425 $D=0
M548 VSS WL<27> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=18960 $D=0
M549 VSS WL<26> 357 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=20495 $D=0
M550 VSS WL<25> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=22030 $D=0
M551 VSS WL<24> 358 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=23565 $D=0
M552 VSS WL<23> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=25100 $D=0
M553 VSS WL<22> 359 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=26635 $D=0
M554 VSS WL<21> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=28170 $D=0
M555 VSS WL<20> 360 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=29705 $D=0
M556 VSS WL<19> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=31240 $D=0
M557 VSS WL<18> 361 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=32775 $D=0
M558 VSS WL<17> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=34310 $D=0
M559 VSS WL<16> 362 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=35845 $D=0
M560 VSS WL<15> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=37800 $D=0
M561 VSS WL<14> 363 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=39335 $D=0
M562 VSS WL<13> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=40870 $D=0
M563 VSS WL<12> 364 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=42405 $D=0
M564 VSS WL<11> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=43940 $D=0
M565 VSS WL<10> 365 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=45475 $D=0
M566 VSS WL<9> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=47010 $D=0
M567 VSS WL<8> 366 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=48545 $D=0
M568 VSS WL<7> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=50080 $D=0
M569 VSS WL<6> 367 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=51615 $D=0
M570 VSS WL<5> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=53150 $D=0
M571 VSS WL<4> 368 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=54685 $D=0
M572 VSS WL<3> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=56220 $D=0
M573 VSS WL<2> 369 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=57755 $D=0
M574 VSS WL<1> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=59290 $D=0
M575 VSS WL<0> 370 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=32685 $Y=60825 $D=0
M576 371 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-37140 $D=0
M577 BL<9> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-35605 $D=0
M578 372 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-34070 $D=0
M579 BL<9> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-32535 $D=0
M580 373 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-31000 $D=0
M581 BL<9> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-29465 $D=0
M582 374 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-27930 $D=0
M583 BL<9> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-26395 $D=0
M584 375 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-24860 $D=0
M585 BL<9> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-23325 $D=0
M586 376 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-21790 $D=0
M587 BL<9> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-20255 $D=0
M588 377 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-18720 $D=0
M589 BL<9> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-17185 $D=0
M590 378 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-15650 $D=0
M591 BL<9> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-14115 $D=0
M592 379 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-12160 $D=0
M593 BL<9> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-10625 $D=0
M594 380 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-9090 $D=0
M595 BL<9> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-7555 $D=0
M596 381 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-6020 $D=0
M597 BL<9> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-4485 $D=0
M598 382 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-2950 $D=0
M599 BL<9> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=-1415 $D=0
M600 383 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=120 $D=0
M601 BL<9> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=1655 $D=0
M602 384 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=3190 $D=0
M603 BL<9> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=4725 $D=0
M604 385 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=6260 $D=0
M605 BL<9> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=7795 $D=0
M606 386 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=9330 $D=0
M607 BL<9> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=10865 $D=0
M608 387 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=12820 $D=0
M609 BL<9> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=14355 $D=0
M610 388 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=15890 $D=0
M611 BL<9> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=17425 $D=0
M612 389 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=18960 $D=0
M613 BL<9> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=20495 $D=0
M614 390 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=22030 $D=0
M615 BL<9> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=23565 $D=0
M616 391 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=25100 $D=0
M617 BL<9> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=26635 $D=0
M618 392 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=28170 $D=0
M619 BL<9> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=29705 $D=0
M620 393 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=31240 $D=0
M621 BL<9> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=32775 $D=0
M622 394 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=34310 $D=0
M623 BL<9> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=35845 $D=0
M624 395 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=37800 $D=0
M625 BL<9> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=39335 $D=0
M626 396 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=40870 $D=0
M627 BL<9> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=42405 $D=0
M628 397 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=43940 $D=0
M629 BL<9> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=45475 $D=0
M630 398 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=47010 $D=0
M631 BL<9> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=48545 $D=0
M632 399 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=50080 $D=0
M633 BL<9> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=51615 $D=0
M634 400 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=53150 $D=0
M635 BL<9> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=54685 $D=0
M636 401 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=56220 $D=0
M637 BL<9> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=57755 $D=0
M638 402 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=59290 $D=0
M639 BL<9> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=33375 $Y=60825 $D=0
M640 VSS WL<63> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-37140 $D=0
M641 VSS WL<62> 403 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-35605 $D=0
M642 VSS WL<61> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-34070 $D=0
M643 VSS WL<60> 404 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-32535 $D=0
M644 VSS WL<59> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-31000 $D=0
M645 VSS WL<58> 405 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-29465 $D=0
M646 VSS WL<57> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-27930 $D=0
M647 VSS WL<56> 406 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-26395 $D=0
M648 VSS WL<55> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-24860 $D=0
M649 VSS WL<54> 407 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-23325 $D=0
M650 VSS WL<53> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-21790 $D=0
M651 VSS WL<52> 408 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-20255 $D=0
M652 VSS WL<51> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-18720 $D=0
M653 VSS WL<50> 409 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-17185 $D=0
M654 VSS WL<49> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-15650 $D=0
M655 VSS WL<48> 410 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-14115 $D=0
M656 VSS WL<47> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-12160 $D=0
M657 VSS WL<46> 411 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-10625 $D=0
M658 VSS WL<45> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-9090 $D=0
M659 VSS WL<44> 412 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-7555 $D=0
M660 VSS WL<43> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-6020 $D=0
M661 VSS WL<42> 413 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-4485 $D=0
M662 VSS WL<41> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-2950 $D=0
M663 VSS WL<40> 414 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=-1415 $D=0
M664 VSS WL<39> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=120 $D=0
M665 VSS WL<38> 415 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=1655 $D=0
M666 VSS WL<37> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=3190 $D=0
M667 VSS WL<36> 416 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=4725 $D=0
M668 VSS WL<35> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=6260 $D=0
M669 VSS WL<34> 417 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=7795 $D=0
M670 VSS WL<33> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=9330 $D=0
M671 VSS WL<32> 418 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=10865 $D=0
M672 VSS WL<31> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=12820 $D=0
M673 VSS WL<30> 419 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=14355 $D=0
M674 VSS WL<29> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=15890 $D=0
M675 VSS WL<28> 420 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=17425 $D=0
M676 VSS WL<27> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=18960 $D=0
M677 VSS WL<26> 421 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=20495 $D=0
M678 VSS WL<25> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=22030 $D=0
M679 VSS WL<24> 422 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=23565 $D=0
M680 VSS WL<23> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=25100 $D=0
M681 VSS WL<22> 423 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=26635 $D=0
M682 VSS WL<21> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=28170 $D=0
M683 VSS WL<20> 424 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=29705 $D=0
M684 VSS WL<19> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=31240 $D=0
M685 VSS WL<18> 425 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=32775 $D=0
M686 VSS WL<17> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=34310 $D=0
M687 VSS WL<16> 426 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=35845 $D=0
M688 VSS WL<15> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=37800 $D=0
M689 VSS WL<14> 427 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=39335 $D=0
M690 VSS WL<13> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=40870 $D=0
M691 VSS WL<12> 428 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=42405 $D=0
M692 VSS WL<11> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=43940 $D=0
M693 VSS WL<10> 429 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=45475 $D=0
M694 VSS WL<9> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=47010 $D=0
M695 VSS WL<8> 430 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=48545 $D=0
M696 VSS WL<7> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=50080 $D=0
M697 VSS WL<6> 431 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=51615 $D=0
M698 VSS WL<5> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=53150 $D=0
M699 VSS WL<4> 432 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=54685 $D=0
M700 VSS WL<3> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=56220 $D=0
M701 VSS WL<2> 433 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=57755 $D=0
M702 VSS WL<1> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=59290 $D=0
M703 VSS WL<0> 434 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=34835 $Y=60825 $D=0
M704 435 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-37140 $D=0
M705 BL<11> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-35605 $D=0
M706 436 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-34070 $D=0
M707 BL<11> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-32535 $D=0
M708 437 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-31000 $D=0
M709 BL<11> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-29465 $D=0
M710 438 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-27930 $D=0
M711 BL<11> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-26395 $D=0
M712 439 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-24860 $D=0
M713 BL<11> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-23325 $D=0
M714 440 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-21790 $D=0
M715 BL<11> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-20255 $D=0
M716 441 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-18720 $D=0
M717 BL<11> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-17185 $D=0
M718 442 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-15650 $D=0
M719 BL<11> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-14115 $D=0
M720 443 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-12160 $D=0
M721 BL<11> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-10625 $D=0
M722 444 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-9090 $D=0
M723 BL<11> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-7555 $D=0
M724 445 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-6020 $D=0
M725 BL<11> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-4485 $D=0
M726 446 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-2950 $D=0
M727 BL<11> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=-1415 $D=0
M728 447 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=120 $D=0
M729 BL<11> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=1655 $D=0
M730 448 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=3190 $D=0
M731 BL<11> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=4725 $D=0
M732 449 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=6260 $D=0
M733 BL<11> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=7795 $D=0
M734 450 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=9330 $D=0
M735 BL<11> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=10865 $D=0
M736 451 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=12820 $D=0
M737 BL<11> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=14355 $D=0
M738 452 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=15890 $D=0
M739 BL<11> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=17425 $D=0
M740 453 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=18960 $D=0
M741 BL<11> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=20495 $D=0
M742 454 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=22030 $D=0
M743 BL<11> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=23565 $D=0
M744 455 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=25100 $D=0
M745 BL<11> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=26635 $D=0
M746 456 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=28170 $D=0
M747 BL<11> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=29705 $D=0
M748 457 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=31240 $D=0
M749 BL<11> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=32775 $D=0
M750 458 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=34310 $D=0
M751 BL<11> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=35845 $D=0
M752 459 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=37800 $D=0
M753 BL<11> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=39335 $D=0
M754 460 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=40870 $D=0
M755 BL<11> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=42405 $D=0
M756 461 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=43940 $D=0
M757 BL<11> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=45475 $D=0
M758 462 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=47010 $D=0
M759 BL<11> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=48545 $D=0
M760 463 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=50080 $D=0
M761 BL<11> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=51615 $D=0
M762 464 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=53150 $D=0
M763 BL<11> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=54685 $D=0
M764 465 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=56220 $D=0
M765 BL<11> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=57755 $D=0
M766 466 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=59290 $D=0
M767 BL<11> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=35525 $Y=60825 $D=0
M768 VSS WL<63> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-37140 $D=0
M769 VSS WL<62> 467 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-35605 $D=0
M770 VSS WL<61> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-34070 $D=0
M771 VSS WL<60> 468 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-32535 $D=0
M772 VSS WL<59> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-31000 $D=0
M773 VSS WL<58> 469 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-29465 $D=0
M774 VSS WL<57> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-27930 $D=0
M775 VSS WL<56> 470 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-26395 $D=0
M776 VSS WL<55> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-24860 $D=0
M777 VSS WL<54> 471 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-23325 $D=0
M778 VSS WL<53> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-21790 $D=0
M779 VSS WL<52> 472 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-20255 $D=0
M780 VSS WL<51> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-18720 $D=0
M781 VSS WL<50> 473 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-17185 $D=0
M782 VSS WL<49> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-15650 $D=0
M783 VSS WL<48> 474 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-14115 $D=0
M784 VSS WL<47> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-12160 $D=0
M785 VSS WL<46> 475 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-10625 $D=0
M786 VSS WL<45> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-9090 $D=0
M787 VSS WL<44> 476 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-7555 $D=0
M788 VSS WL<43> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-6020 $D=0
M789 VSS WL<42> 477 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-4485 $D=0
M790 VSS WL<41> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-2950 $D=0
M791 VSS WL<40> 478 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=-1415 $D=0
M792 VSS WL<39> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=120 $D=0
M793 VSS WL<38> 479 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=1655 $D=0
M794 VSS WL<37> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=3190 $D=0
M795 VSS WL<36> 480 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=4725 $D=0
M796 VSS WL<35> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=6260 $D=0
M797 VSS WL<34> 481 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=7795 $D=0
M798 VSS WL<33> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=9330 $D=0
M799 VSS WL<32> 482 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=10865 $D=0
M800 VSS WL<31> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=12820 $D=0
M801 VSS WL<30> 483 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=14355 $D=0
M802 VSS WL<29> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=15890 $D=0
M803 VSS WL<28> 484 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=17425 $D=0
M804 VSS WL<27> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=18960 $D=0
M805 VSS WL<26> 485 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=20495 $D=0
M806 VSS WL<25> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=22030 $D=0
M807 VSS WL<24> 486 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=23565 $D=0
M808 VSS WL<23> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=25100 $D=0
M809 VSS WL<22> 487 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=26635 $D=0
M810 VSS WL<21> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=28170 $D=0
M811 VSS WL<20> 488 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=29705 $D=0
M812 VSS WL<19> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=31240 $D=0
M813 VSS WL<18> 489 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=32775 $D=0
M814 VSS WL<17> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=34310 $D=0
M815 VSS WL<16> 490 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=35845 $D=0
M816 VSS WL<15> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=37800 $D=0
M817 VSS WL<14> 491 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=39335 $D=0
M818 VSS WL<13> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=40870 $D=0
M819 VSS WL<12> 492 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=42405 $D=0
M820 VSS WL<11> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=43940 $D=0
M821 VSS WL<10> 493 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=45475 $D=0
M822 VSS WL<9> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=47010 $D=0
M823 VSS WL<8> 494 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=48545 $D=0
M824 VSS WL<7> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=50080 $D=0
M825 VSS WL<6> 495 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=51615 $D=0
M826 VSS WL<5> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=53150 $D=0
M827 VSS WL<4> 496 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=54685 $D=0
M828 VSS WL<3> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=56220 $D=0
M829 VSS WL<2> 497 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=57755 $D=0
M830 VSS WL<1> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=59290 $D=0
M831 VSS WL<0> 498 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=36985 $Y=60825 $D=0
M832 499 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-37140 $D=0
M833 BL<13> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-35605 $D=0
M834 500 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-34070 $D=0
M835 BL<13> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-32535 $D=0
M836 501 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-31000 $D=0
M837 BL<13> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-29465 $D=0
M838 502 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-27930 $D=0
M839 BL<13> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-26395 $D=0
M840 503 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-24860 $D=0
M841 BL<13> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-23325 $D=0
M842 504 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-21790 $D=0
M843 BL<13> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-20255 $D=0
M844 505 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-18720 $D=0
M845 BL<13> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-17185 $D=0
M846 506 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-15650 $D=0
M847 BL<13> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-14115 $D=0
M848 507 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-12160 $D=0
M849 BL<13> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-10625 $D=0
M850 508 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-9090 $D=0
M851 BL<13> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-7555 $D=0
M852 509 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-6020 $D=0
M853 BL<13> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-4485 $D=0
M854 510 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-2950 $D=0
M855 BL<13> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=-1415 $D=0
M856 511 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=120 $D=0
M857 BL<13> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=1655 $D=0
M858 512 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=3190 $D=0
M859 BL<13> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=4725 $D=0
M860 513 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=6260 $D=0
M861 BL<13> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=7795 $D=0
M862 514 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=9330 $D=0
M863 BL<13> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=10865 $D=0
M864 515 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=12820 $D=0
M865 BL<13> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=14355 $D=0
M866 516 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=15890 $D=0
M867 BL<13> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=17425 $D=0
M868 517 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=18960 $D=0
M869 BL<13> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=20495 $D=0
M870 518 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=22030 $D=0
M871 BL<13> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=23565 $D=0
M872 519 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=25100 $D=0
M873 BL<13> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=26635 $D=0
M874 520 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=28170 $D=0
M875 BL<13> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=29705 $D=0
M876 521 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=31240 $D=0
M877 BL<13> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=32775 $D=0
M878 522 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=34310 $D=0
M879 BL<13> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=35845 $D=0
M880 523 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=37800 $D=0
M881 BL<13> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=39335 $D=0
M882 524 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=40870 $D=0
M883 BL<13> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=42405 $D=0
M884 525 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=43940 $D=0
M885 BL<13> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=45475 $D=0
M886 526 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=47010 $D=0
M887 BL<13> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=48545 $D=0
M888 527 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=50080 $D=0
M889 BL<13> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=51615 $D=0
M890 528 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=53150 $D=0
M891 BL<13> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=54685 $D=0
M892 529 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=56220 $D=0
M893 BL<13> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=57755 $D=0
M894 530 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=59290 $D=0
M895 BL<13> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=37675 $Y=60825 $D=0
M896 VSS WL<63> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-37140 $D=0
M897 VSS WL<62> 531 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-35605 $D=0
M898 VSS WL<61> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-34070 $D=0
M899 VSS WL<60> 532 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-32535 $D=0
M900 VSS WL<59> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-31000 $D=0
M901 VSS WL<58> 533 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-29465 $D=0
M902 VSS WL<57> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-27930 $D=0
M903 VSS WL<56> 534 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-26395 $D=0
M904 VSS WL<55> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-24860 $D=0
M905 VSS WL<54> 535 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-23325 $D=0
M906 VSS WL<53> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-21790 $D=0
M907 VSS WL<52> 536 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-20255 $D=0
M908 VSS WL<51> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-18720 $D=0
M909 VSS WL<50> 537 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-17185 $D=0
M910 VSS WL<49> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-15650 $D=0
M911 VSS WL<48> 538 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-14115 $D=0
M912 VSS WL<47> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-12160 $D=0
M913 VSS WL<46> 539 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-10625 $D=0
M914 VSS WL<45> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-9090 $D=0
M915 VSS WL<44> 540 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-7555 $D=0
M916 VSS WL<43> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-6020 $D=0
M917 VSS WL<42> 541 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-4485 $D=0
M918 VSS WL<41> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-2950 $D=0
M919 VSS WL<40> 542 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=-1415 $D=0
M920 VSS WL<39> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=120 $D=0
M921 VSS WL<38> 543 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=1655 $D=0
M922 VSS WL<37> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=3190 $D=0
M923 VSS WL<36> 544 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=4725 $D=0
M924 VSS WL<35> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=6260 $D=0
M925 VSS WL<34> 545 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=7795 $D=0
M926 VSS WL<33> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=9330 $D=0
M927 VSS WL<32> 546 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=10865 $D=0
M928 VSS WL<31> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=12820 $D=0
M929 VSS WL<30> 547 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=14355 $D=0
M930 VSS WL<29> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=15890 $D=0
M931 VSS WL<28> 548 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=17425 $D=0
M932 VSS WL<27> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=18960 $D=0
M933 VSS WL<26> 549 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=20495 $D=0
M934 VSS WL<25> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=22030 $D=0
M935 VSS WL<24> 550 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=23565 $D=0
M936 VSS WL<23> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=25100 $D=0
M937 VSS WL<22> 551 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=26635 $D=0
M938 VSS WL<21> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=28170 $D=0
M939 VSS WL<20> 552 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=29705 $D=0
M940 VSS WL<19> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=31240 $D=0
M941 VSS WL<18> 553 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=32775 $D=0
M942 VSS WL<17> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=34310 $D=0
M943 VSS WL<16> 554 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=35845 $D=0
M944 VSS WL<15> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=37800 $D=0
M945 VSS WL<14> 555 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=39335 $D=0
M946 VSS WL<13> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=40870 $D=0
M947 VSS WL<12> 556 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=42405 $D=0
M948 VSS WL<11> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=43940 $D=0
M949 VSS WL<10> 557 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=45475 $D=0
M950 VSS WL<9> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=47010 $D=0
M951 VSS WL<8> 558 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=48545 $D=0
M952 VSS WL<7> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=50080 $D=0
M953 VSS WL<6> 559 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=51615 $D=0
M954 VSS WL<5> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=53150 $D=0
M955 VSS WL<4> 560 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=54685 $D=0
M956 VSS WL<3> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=56220 $D=0
M957 VSS WL<2> 561 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=57755 $D=0
M958 VSS WL<1> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=59290 $D=0
M959 VSS WL<0> 562 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=39135 $Y=60825 $D=0
M960 564 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-37140 $D=0
M961 BL<15> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-35605 $D=0
M962 565 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-34070 $D=0
M963 BL<15> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-32535 $D=0
M964 566 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-31000 $D=0
M965 BL<15> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-29465 $D=0
M966 567 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-27930 $D=0
M967 BL<15> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-26395 $D=0
M968 568 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-24860 $D=0
M969 BL<15> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-23325 $D=0
M970 569 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-21790 $D=0
M971 BL<15> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-20255 $D=0
M972 570 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-18720 $D=0
M973 BL<15> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-17185 $D=0
M974 571 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-15650 $D=0
M975 BL<15> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-14115 $D=0
M976 572 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-12160 $D=0
M977 BL<15> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-10625 $D=0
M978 573 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-9090 $D=0
M979 BL<15> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-7555 $D=0
M980 574 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-6020 $D=0
M981 BL<15> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-4485 $D=0
M982 575 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-2950 $D=0
M983 BL<15> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=-1415 $D=0
M984 576 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=120 $D=0
M985 BL<15> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=1655 $D=0
M986 577 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=3190 $D=0
M987 BL<15> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=4725 $D=0
M988 578 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=6260 $D=0
M989 BL<15> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=7795 $D=0
M990 579 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=9330 $D=0
M991 BL<15> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=10865 $D=0
M992 580 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=12820 $D=0
M993 BL<15> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=14355 $D=0
M994 581 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=15890 $D=0
M995 BL<15> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=17425 $D=0
M996 582 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=18960 $D=0
M997 BL<15> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=20495 $D=0
M998 583 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=22030 $D=0
M999 BL<15> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=23565 $D=0
M1000 584 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=25100 $D=0
M1001 BL<15> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=26635 $D=0
M1002 585 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=28170 $D=0
M1003 BL<15> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=29705 $D=0
M1004 586 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=31240 $D=0
M1005 BL<15> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=32775 $D=0
M1006 587 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=34310 $D=0
M1007 BL<15> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=35845 $D=0
M1008 588 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=37800 $D=0
M1009 BL<15> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=39335 $D=0
M1010 589 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=40870 $D=0
M1011 BL<15> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=42405 $D=0
M1012 590 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=43940 $D=0
M1013 BL<15> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=45475 $D=0
M1014 591 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=47010 $D=0
M1015 BL<15> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=48545 $D=0
M1016 592 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=50080 $D=0
M1017 BL<15> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=51615 $D=0
M1018 593 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=53150 $D=0
M1019 BL<15> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=54685 $D=0
M1020 594 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=56220 $D=0
M1021 BL<15> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=57755 $D=0
M1022 595 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=59290 $D=0
M1023 BL<15> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=39825 $Y=60825 $D=0
M1024 VDD pre_b BL<0> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=24085 $Y=-40540 $D=1
M1025 BL<1> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=24775 $Y=-40540 $D=1
M1026 VDD pre_b BL<2> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=26235 $Y=-40540 $D=1
M1027 BL<3> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=26925 $Y=-40540 $D=1
M1028 VDD pre_b BL<4> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=28385 $Y=-40540 $D=1
M1029 BL<5> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=29075 $Y=-40540 $D=1
M1030 VDD pre_b BL<6> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=30535 $Y=-40540 $D=1
M1031 BL<7> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=31225 $Y=-40540 $D=1
M1032 VDD pre_b BL<8> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=32685 $Y=-40540 $D=1
M1033 BL<9> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=33375 $Y=-40540 $D=1
M1034 VDD pre_b BL<10> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=34835 $Y=-40540 $D=1
M1035 BL<11> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=35525 $Y=-40540 $D=1
M1036 VDD pre_b BL<12> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=36985 $Y=-40540 $D=1
M1037 BL<13> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=37675 $Y=-40540 $D=1
M1038 VDD pre_b BL<14> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=39135 $Y=-40540 $D=1
M1039 BL<15> pre_b VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=39825 $Y=-40540 $D=1
.ENDS
***************************************
