* File: hw3_part1.pex.spi
* Created: Tue Nov 23 22:04:25 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw3_part1.pex.spi.pex"
.subckt hw3_part1  Q VSS VDD QB CLK R S
* 
* S	S
* R	R
* CLK	CLK
* QB	QB
* VDD	VDD
* VSS	VSS
* Q	Q
MM0 N_Q_MM0_d N_QB_MM0_g N_VDD_MM0_s N_VDD_MM0_b P_18 L=1.8e-07 W=2e-06
+ AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06
MM3 N_QB_MM3_d N_Q_MM3_g N_VDD_MM3_s N_VDD_MM0_b P_18 L=1.8e-07 W=2e-06
+ AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06
MM1 N_Q_MM1_d N_QB_MM1_g N_VSS_MM1_s N_VSS_MM1_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM2 N_QB_MM2_d N_Q_MM2_g N_VSS_MM2_s N_VSS_MM1_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM4 N_R_MM4_d N_CLK_MM4_g N_QB_MM4_s N_VSS_MM1_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM5 N_S_MM5_d N_CLK_MM5_g N_Q_MM5_s N_VSS_MM1_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
*
.include "hw3_part1.pex.spi.HW3_PART1.pxi"
*
.ends
*
*
