* SPICE NETLIST
***************************************

*.CALIBRE ABORT_INFO SOFTCHK
.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT mos_unit2
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT mos_unit
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Final_SA 1 2 3 4 5 6 7
** N=10 EP=7 IP=40 FDC=12
M0 9 4 8 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-2175 $Y=-410 $D=0
M1 5 3 8 5 N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-1310 $Y=-1590 $D=0
M2 2 1 9 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-715 $Y=-410 $D=0
M3 8 3 5 5 N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-620 $Y=-1590 $D=0
M4 5 3 8 5 N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=70 $Y=-1590 $D=0
M5 10 2 1 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=745 $Y=-410 $D=0
M6 8 3 5 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=760 $Y=-1590 $D=0
M7 8 6 10 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=2205 $Y=-410 $D=0
M8 2 3 7 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-2175 $Y=1410 $D=1
M9 2 1 7 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-715 $Y=1410 $D=1
M10 7 2 1 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=745 $Y=1410 $D=1
M11 7 3 1 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=2205 $Y=1410 $D=1
.ENDS
***************************************
.SUBCKT final_mos_unit
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT inv_final 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 2 2 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-65 $Y=-2195 $D=0
M1 4 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-65 $Y=-490 $D=1
.ENDS
***************************************
.SUBCKT final_and 1 2 3 4 5
** N=7 EP=5 IP=28 FDC=6
M0 7 2 4 4 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=8825 $Y=670 $D=0
M1 6 1 7 4 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=8825 $Y=2130 $D=0
M2 6 2 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10465 $Y=670 $D=1
M3 6 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10465 $Y=2130 $D=1
X12 6 4 3 5 inv_final $T=14700 2115 0 0 $X=13540 $Y=-1150
.ENDS
***************************************
.SUBCKT inv_1u5_0u5 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 2 2 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-65 $Y=-2195 $D=0
M1 4 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-65 $Y=-490 $D=1
.ENDS
***************************************
.SUBCKT ICV_1
** N=6 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT nand4_final
** N=9 EP=0 IP=24 FDC=0
.ENDS
***************************************
.SUBCKT Ydecoder_final 1 2 3 4 5 6 7 8 9 10 11 12 13
** N=40 EP=13 IP=84 FDC=70
M0 17 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=-1665 $D=0
M1 21 3 17 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=-205 $D=0
M2 25 2 21 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=1255 $D=0
M3 4 14 25 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=2715 $D=0
M4 18 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=4355 $D=0
M5 22 16 18 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=5815 $D=0
M6 26 2 22 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=7275 $D=0
M7 5 14 26 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=8735 $D=0
M8 19 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=10375 $D=0
M9 23 3 19 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=11835 $D=0
M10 27 15 23 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=13295 $D=0
M11 6 14 27 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=14755 $D=0
M12 20 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=16395 $D=0
M13 24 16 20 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=17855 $D=0
M14 28 15 24 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=19315 $D=0
M15 7 14 28 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=20775 $D=0
M16 29 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=-1645 $D=0
M17 33 3 29 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=-185 $D=0
M18 37 2 33 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=1275 $D=0
M19 8 1 37 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=2735 $D=0
M20 30 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=4375 $D=0
M21 34 16 30 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=5835 $D=0
M22 38 2 34 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=7295 $D=0
M23 9 1 38 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=8755 $D=0
M24 31 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=10395 $D=0
M25 35 3 31 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=11855 $D=0
M26 39 15 35 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=13315 $D=0
M27 10 1 39 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=14775 $D=0
M28 32 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=16415 $D=0
M29 36 16 32 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=17875 $D=0
M30 40 15 36 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=19335 $D=0
M31 11 1 40 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=20795 $D=0
M32 4 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=-1665 $D=1
M33 4 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=-205 $D=1
M34 4 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=1255 $D=1
M35 4 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=2715 $D=1
M36 5 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=4355 $D=1
M37 5 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=5815 $D=1
M38 5 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=7275 $D=1
M39 5 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=8735 $D=1
M40 6 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=10375 $D=1
M41 6 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=11835 $D=1
M42 6 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=13295 $D=1
M43 6 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=14755 $D=1
M44 7 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=16395 $D=1
M45 7 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=17855 $D=1
M46 7 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=19315 $D=1
M47 7 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=20775 $D=1
M48 8 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=-1645 $D=1
M49 8 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=-185 $D=1
M50 8 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=1275 $D=1
M51 8 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=2735 $D=1
M52 9 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=4375 $D=1
M53 9 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=5835 $D=1
M54 9 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=7295 $D=1
M55 9 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=8755 $D=1
M56 10 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=10395 $D=1
M57 10 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=11855 $D=1
M58 10 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=13315 $D=1
M59 10 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=14775 $D=1
M60 11 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=16415 $D=1
M61 11 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=17875 $D=1
M62 11 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=19335 $D=1
M63 11 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=20795 $D=1
X64 3 13 12 16 inv_1u5_0u5 $T=985 1015 0 0 $X=-175 $Y=-2250
X65 2 13 12 15 inv_1u5_0u5 $T=985 7265 0 0 $X=-175 $Y=4000
X66 1 13 12 14 inv_1u5_0u5 $T=985 19305 0 0 $X=-175 $Y=16040
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X0 1 2 3 4 inv_final $T=0 0 0 0 $X=-1160 $Y=-3265
X1 4 2 3 5 inv_final $T=1600 0 0 0 $X=440 $Y=-3265
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5
** N=7 EP=5 IP=10 FDC=8
X0 1 2 3 6 7 ICV_2 $T=0 0 0 0 $X=-1160 $Y=-3265
X1 7 2 3 4 5 ICV_2 $T=3200 0 0 0 $X=2040 $Y=-3265
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4
** N=7 EP=4 IP=10 FDC=16
X0 1 2 3 5 6 ICV_3 $T=0 0 0 0 $X=-1160 $Y=-3265
X1 6 2 3 7 4 ICV_3 $T=6400 0 0 0 $X=5240 $Y=-3265
.ENDS
***************************************
.SUBCKT FInal_FF 1 2 3 4 5 6
** N=15 EP=6 IP=16 FDC=20
M0 9 1 7 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-2285 $Y=-2400 $D=0
M1 11 2 3 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=1670 $Y=-2400 $D=0
M2 7 12 11 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=3170 $Y=-2400 $D=0
M3 8 2 12 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=5540 $Y=-1425 $D=0
M4 13 1 3 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=9425 $Y=-2400 $D=0
M5 8 15 13 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10925 $Y=-2400 $D=0
M6 9 2 7 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-2285 $Y=-5120 $D=1
M7 10 1 4 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=1570 $Y=-5120 $D=1
M8 7 12 10 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=3170 $Y=-5120 $D=1
M9 8 1 12 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=5540 $Y=295 $D=1
M10 14 2 4 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=9425 $Y=-5120 $D=1
M11 8 15 14 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=10925 $Y=-5120 $D=1
X12 5 3 4 9 inv_1u5_0u5 $T=-2220 1570 0 0 $X=-3380 $Y=-1695
X13 7 3 4 12 inv_1u5_0u5 $T=1735 1565 0 0 $X=575 $Y=-1700
X14 8 3 4 15 inv_1u5_0u5 $T=9490 1565 0 0 $X=8330 $Y=-1700
X15 15 3 4 6 inv_1u5_0u5 $T=13725 1565 0 0 $X=12565 $Y=-1700
.ENDS
***************************************
.SUBCKT Final_all_v1 YOUT<0> YOUT<1> YOUT<2> YOUT<3> YOUT<4> YOUT<5> YOUT<6> YOUT<7> Dout<0> SO<0> Dout<1> SO<1> VDD CLK WL_EN SAEN BL<0> BL<1> BL<2> BL<3>
+ BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15> VSS X_sel<5> X_sel<2> X_sel<4> X_sel<1> X_sel<3> X_sel<0> WL<63>
+ WL<62> WL<61> WL<60> WL<59> WL<58> WL<57> WL<56> WL<55> WL<54> WL<53> WL<52> WL<51> WL<50> WL<49> WL<48> WL<47> WL<46> WL<45> WL<44> WL<43>
+ WL<42> WL<41> WL<40> WL<39> WL<38> WL<37> WL<36> WL<35> WL<34> WL<33> WL<32> WL<31> WL<30> WL<29> WL<28> WL<27> WL<26> WL<25> WL<24> WL<23>
+ WL<22> WL<21> WL<20> WL<19> WL<18> WL<17> WL<16> WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3>
+ WL<2> WL<1> WL<0> DL<0> DL<1> Y_sel<0> Y_sel<2> Y_sel<1> Vref A<2> A<1> A<0> A<6> A<7> A<8> A<3> A<4> A<5>
** N=811 EP=118 IP=139 FDC=1897
D0 VSS VDD DN AREA=5.64e-13 PJ=3.34e-06 $X=-25674 $Y=-31450 $D=31
M1 83 X_sel<3> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=7260 $D=0
M2 81 X_sel<4> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=19300 $D=0
M3 85 X_sel<5> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=31340 $D=0
M4 84 X_sel<0> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=55940 $D=0
M5 82 X_sel<1> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=67980 $D=0
M6 86 X_sel<2> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=80020 $D=0
M7 168 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-11510 $D=0
M8 169 X_sel<3> 168 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-10050 $D=0
M9 170 X_sel<4> 169 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-8590 $D=0
M10 16 X_sel<5> 170 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-7130 $D=0
M11 171 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-5490 $D=0
M12 172 83 171 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-4030 $D=0
M13 173 X_sel<4> 172 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-2570 $D=0
M14 17 X_sel<5> 173 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-1110 $D=0
M15 174 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=530 $D=0
M16 175 X_sel<3> 174 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=1990 $D=0
M17 176 81 175 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=3450 $D=0
M18 18 X_sel<5> 176 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=4910 $D=0
M19 177 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=6550 $D=0
M20 178 83 177 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=8010 $D=0
M21 179 81 178 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=9470 $D=0
M22 19 X_sel<5> 179 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=10930 $D=0
M23 180 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=12570 $D=0
M24 181 X_sel<3> 180 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=14030 $D=0
M25 182 X_sel<4> 181 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=15490 $D=0
M26 20 85 182 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=16950 $D=0
M27 183 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=18590 $D=0
M28 184 83 183 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=20050 $D=0
M29 185 X_sel<4> 184 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=21510 $D=0
M30 21 85 185 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=22970 $D=0
M31 186 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=24610 $D=0
M32 187 X_sel<3> 186 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=26070 $D=0
M33 188 81 187 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=27530 $D=0
M34 22 85 188 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=28990 $D=0
M35 189 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=30630 $D=0
M36 190 83 189 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=32090 $D=0
M37 191 81 190 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=33550 $D=0
M38 23 85 191 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=35010 $D=0
M39 192 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=37170 $D=0
M40 193 X_sel<0> 192 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=38630 $D=0
M41 194 X_sel<1> 193 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=40090 $D=0
M42 24 X_sel<2> 194 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=41550 $D=0
M43 195 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=43190 $D=0
M44 196 84 195 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=44650 $D=0
M45 197 X_sel<1> 196 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=46110 $D=0
M46 25 X_sel<2> 197 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=47570 $D=0
M47 198 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=49210 $D=0
M48 199 X_sel<0> 198 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=50670 $D=0
M49 200 82 199 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=52130 $D=0
M50 26 X_sel<2> 200 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=53590 $D=0
M51 201 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=55230 $D=0
M52 202 84 201 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=56690 $D=0
M53 203 82 202 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=58150 $D=0
M54 27 X_sel<2> 203 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=59610 $D=0
M55 204 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=61250 $D=0
M56 205 X_sel<0> 204 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=62710 $D=0
M57 206 X_sel<1> 205 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=64170 $D=0
M58 28 86 206 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=65630 $D=0
M59 207 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=67270 $D=0
M60 208 84 207 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=68730 $D=0
M61 209 X_sel<1> 208 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=70190 $D=0
M62 29 86 209 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=71650 $D=0
M63 210 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=73290 $D=0
M64 211 X_sel<0> 210 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=74750 $D=0
M65 212 82 211 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=76210 $D=0
M66 30 86 212 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=77670 $D=0
M67 213 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=79310 $D=0
M68 214 84 213 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=80770 $D=0
M69 215 82 214 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=82230 $D=0
M70 31 86 215 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=83690 $D=0
M71 WL<63> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-13505 $D=0
M72 WL<62> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-11970 $D=0
M73 WL<61> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-10435 $D=0
M74 WL<60> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-8900 $D=0
M75 WL<59> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-7365 $D=0
M76 WL<58> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-5830 $D=0
M77 WL<57> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-4295 $D=0
M78 WL<56> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-2760 $D=0
M79 WL<55> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-1225 $D=0
M80 WL<54> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=310 $D=0
M81 WL<53> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=1845 $D=0
M82 WL<52> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=3380 $D=0
M83 WL<51> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=4915 $D=0
M84 WL<50> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=6450 $D=0
M85 WL<49> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=7985 $D=0
M86 WL<48> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=9520 $D=0
M87 WL<47> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=11475 $D=0
M88 WL<46> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=13010 $D=0
M89 WL<45> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=14545 $D=0
M90 WL<44> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=16080 $D=0
M91 WL<43> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=17615 $D=0
M92 WL<42> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=19150 $D=0
M93 WL<41> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=20685 $D=0
M94 WL<40> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=22220 $D=0
M95 WL<39> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=23755 $D=0
M96 WL<38> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=25290 $D=0
M97 WL<37> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=26825 $D=0
M98 WL<36> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=28360 $D=0
M99 WL<35> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=29895 $D=0
M100 WL<34> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=31430 $D=0
M101 WL<33> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=32965 $D=0
M102 WL<32> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=34500 $D=0
M103 WL<31> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=36455 $D=0
M104 WL<30> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=37990 $D=0
M105 WL<29> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=39525 $D=0
M106 WL<28> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=41060 $D=0
M107 WL<27> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=42595 $D=0
M108 WL<26> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=44130 $D=0
M109 WL<25> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=45665 $D=0
M110 WL<24> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=47200 $D=0
M111 WL<23> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=48735 $D=0
M112 WL<22> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=50270 $D=0
M113 WL<21> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=51805 $D=0
M114 WL<20> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=53340 $D=0
M115 WL<19> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=54875 $D=0
M116 WL<18> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=56410 $D=0
M117 WL<17> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=57945 $D=0
M118 WL<16> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=59480 $D=0
M119 WL<15> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=61435 $D=0
M120 WL<14> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=62970 $D=0
M121 WL<13> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=64505 $D=0
M122 WL<12> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=66040 $D=0
M123 WL<11> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=67575 $D=0
M124 WL<10> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=69110 $D=0
M125 WL<9> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=70645 $D=0
M126 WL<8> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=72180 $D=0
M127 WL<7> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=73715 $D=0
M128 WL<6> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=75250 $D=0
M129 WL<5> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=76785 $D=0
M130 WL<4> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=78320 $D=0
M131 WL<3> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=79855 $D=0
M132 WL<2> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=81390 $D=0
M133 WL<1> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=82925 $D=0
M134 WL<0> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=84460 $D=0
M135 WL<63> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-13505 $D=0
M136 WL<62> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-11970 $D=0
M137 WL<61> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-10435 $D=0
M138 WL<60> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-8900 $D=0
M139 WL<59> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-7365 $D=0
M140 WL<58> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-5830 $D=0
M141 WL<57> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-4295 $D=0
M142 WL<56> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-2760 $D=0
M143 WL<55> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-1225 $D=0
M144 WL<54> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=310 $D=0
M145 WL<53> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=1845 $D=0
M146 WL<52> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=3380 $D=0
M147 WL<51> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=4915 $D=0
M148 WL<50> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=6450 $D=0
M149 WL<49> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=7985 $D=0
M150 WL<48> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=9520 $D=0
M151 WL<47> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=11475 $D=0
M152 WL<46> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=13010 $D=0
M153 WL<45> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=14545 $D=0
M154 WL<44> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=16080 $D=0
M155 WL<43> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=17615 $D=0
M156 WL<42> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=19150 $D=0
M157 WL<41> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=20685 $D=0
M158 WL<40> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=22220 $D=0
M159 WL<39> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=23755 $D=0
M160 WL<38> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=25290 $D=0
M161 WL<37> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=26825 $D=0
M162 WL<36> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=28360 $D=0
M163 WL<35> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=29895 $D=0
M164 WL<34> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=31430 $D=0
M165 WL<33> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=32965 $D=0
M166 WL<32> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=34500 $D=0
M167 WL<31> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=36455 $D=0
M168 WL<30> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=37990 $D=0
M169 WL<29> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=39525 $D=0
M170 WL<28> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=41060 $D=0
M171 WL<27> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=42595 $D=0
M172 WL<26> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=44130 $D=0
M173 WL<25> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=45665 $D=0
M174 WL<24> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=47200 $D=0
M175 WL<23> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=48735 $D=0
M176 WL<22> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=50270 $D=0
M177 WL<21> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=51805 $D=0
M178 WL<20> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=53340 $D=0
M179 WL<19> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=54875 $D=0
M180 WL<18> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=56410 $D=0
M181 WL<17> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=57945 $D=0
M182 WL<16> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=59480 $D=0
M183 WL<15> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=61435 $D=0
M184 WL<14> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=62970 $D=0
M185 WL<13> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=64505 $D=0
M186 WL<12> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=66040 $D=0
M187 WL<11> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=67575 $D=0
M188 WL<10> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=69110 $D=0
M189 WL<9> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=70645 $D=0
M190 WL<8> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=72180 $D=0
M191 WL<7> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=73715 $D=0
M192 WL<6> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=75250 $D=0
M193 WL<5> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=76785 $D=0
M194 WL<4> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=78320 $D=0
M195 WL<3> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=79855 $D=0
M196 WL<2> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=81390 $D=0
M197 WL<1> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=82925 $D=0
M198 WL<0> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=84460 $D=0
M199 VSS WL<63> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-13645 $D=0
M200 VSS WL<62> 280 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-12110 $D=0
M201 VSS WL<61> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-10575 $D=0
M202 VSS WL<60> 281 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-9040 $D=0
M203 VSS WL<59> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-7505 $D=0
M204 VSS WL<58> 282 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-5970 $D=0
M205 VSS WL<57> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-4435 $D=0
M206 VSS WL<56> 283 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-2900 $D=0
M207 VSS WL<55> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-1365 $D=0
M208 VSS WL<54> 284 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=170 $D=0
M209 VSS WL<53> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=1705 $D=0
M210 VSS WL<52> 285 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=3240 $D=0
M211 VSS WL<51> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=4775 $D=0
M212 VSS WL<50> 286 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=6310 $D=0
M213 VSS WL<49> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=7845 $D=0
M214 VSS WL<48> 287 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=9380 $D=0
M215 VSS WL<47> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=11335 $D=0
M216 VSS WL<46> 288 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=12870 $D=0
M217 VSS WL<45> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=14405 $D=0
M218 VSS WL<44> 289 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=15940 $D=0
M219 VSS WL<43> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=17475 $D=0
M220 VSS WL<42> 290 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=19010 $D=0
M221 VSS WL<41> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=20545 $D=0
M222 VSS WL<40> 291 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=22080 $D=0
M223 VSS WL<39> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=23615 $D=0
M224 VSS WL<38> 292 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=25150 $D=0
M225 VSS WL<37> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=26685 $D=0
M226 VSS WL<36> 293 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=28220 $D=0
M227 VSS WL<35> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=29755 $D=0
M228 VSS WL<34> 294 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=31290 $D=0
M229 VSS WL<33> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=32825 $D=0
M230 VSS WL<32> 295 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=34360 $D=0
M231 VSS WL<31> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=36315 $D=0
M232 VSS WL<30> 296 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=37850 $D=0
M233 VSS WL<29> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=39385 $D=0
M234 VSS WL<28> 297 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=40920 $D=0
M235 VSS WL<27> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=42455 $D=0
M236 VSS WL<26> 298 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=43990 $D=0
M237 VSS WL<25> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=45525 $D=0
M238 VSS WL<24> 299 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=47060 $D=0
M239 VSS WL<23> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=48595 $D=0
M240 VSS WL<22> 300 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=50130 $D=0
M241 VSS WL<21> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=51665 $D=0
M242 VSS WL<20> 301 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=53200 $D=0
M243 VSS WL<19> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=54735 $D=0
M244 VSS WL<18> 302 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=56270 $D=0
M245 VSS WL<17> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=57805 $D=0
M246 VSS WL<16> 303 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=59340 $D=0
M247 VSS WL<15> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=61295 $D=0
M248 VSS WL<14> 304 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=62830 $D=0
M249 VSS WL<13> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=64365 $D=0
M250 VSS WL<12> 305 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=65900 $D=0
M251 VSS WL<11> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=67435 $D=0
M252 VSS WL<10> 306 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=68970 $D=0
M253 VSS WL<9> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=70505 $D=0
M254 VSS WL<8> 307 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=72040 $D=0
M255 VSS WL<7> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=73575 $D=0
M256 VSS WL<6> 308 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=75110 $D=0
M257 VSS WL<5> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=76645 $D=0
M258 VSS WL<4> 309 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=78180 $D=0
M259 VSS WL<3> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=79715 $D=0
M260 VSS WL<2> 310 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=81250 $D=0
M261 VSS WL<1> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=82785 $D=0
M262 VSS WL<0> 311 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=84320 $D=0
M263 36 YOUT<1> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27314 $Y=-35060 $D=0
M264 37 YOUT<0> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27314 $Y=-25360 $D=0
M265 154 36 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27129 $Y=-37026 $D=0
M266 BL<0> 37 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27129 $Y=-27326 $D=0
M267 312 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-13645 $D=0
M268 BL<1> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-12110 $D=0
M269 313 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-10575 $D=0
M270 BL<1> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-9040 $D=0
M271 314 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-7505 $D=0
M272 BL<1> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-5970 $D=0
M273 315 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-4435 $D=0
M274 BL<1> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-2900 $D=0
M275 316 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-1365 $D=0
M276 BL<1> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=170 $D=0
M277 317 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=1705 $D=0
M278 BL<1> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=3240 $D=0
M279 318 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=4775 $D=0
M280 BL<1> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=6310 $D=0
M281 319 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=7845 $D=0
M282 BL<1> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=9380 $D=0
M283 320 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=11335 $D=0
M284 BL<1> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=12870 $D=0
M285 321 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=14405 $D=0
M286 BL<1> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=15940 $D=0
M287 322 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=17475 $D=0
M288 BL<1> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=19010 $D=0
M289 323 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=20545 $D=0
M290 BL<1> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=22080 $D=0
M291 324 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=23615 $D=0
M292 BL<1> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=25150 $D=0
M293 325 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=26685 $D=0
M294 BL<1> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=28220 $D=0
M295 326 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=29755 $D=0
M296 BL<1> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=31290 $D=0
M297 327 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=32825 $D=0
M298 BL<1> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=34360 $D=0
M299 328 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=36315 $D=0
M300 BL<1> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=37850 $D=0
M301 329 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=39385 $D=0
M302 BL<1> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=40920 $D=0
M303 330 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=42455 $D=0
M304 BL<1> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=43990 $D=0
M305 331 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=45525 $D=0
M306 BL<1> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=47060 $D=0
M307 332 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=48595 $D=0
M308 BL<1> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=50130 $D=0
M309 333 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=51665 $D=0
M310 BL<1> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=53200 $D=0
M311 334 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=54735 $D=0
M312 BL<1> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=56270 $D=0
M313 335 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=57805 $D=0
M314 BL<1> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=59340 $D=0
M315 336 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=61295 $D=0
M316 BL<1> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=62830 $D=0
M317 337 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=64365 $D=0
M318 BL<1> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=65900 $D=0
M319 338 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=67435 $D=0
M320 BL<1> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=68970 $D=0
M321 339 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=70505 $D=0
M322 BL<1> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=72040 $D=0
M323 340 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=73575 $D=0
M324 BL<1> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=75110 $D=0
M325 341 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=76645 $D=0
M326 BL<1> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=78180 $D=0
M327 342 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=79715 $D=0
M328 BL<1> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=81250 $D=0
M329 343 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=82785 $D=0
M330 BL<1> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=84320 $D=0
M331 VSS WL<63> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-13645 $D=0
M332 VSS WL<62> 344 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-12110 $D=0
M333 VSS WL<61> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-10575 $D=0
M334 VSS WL<60> 345 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-9040 $D=0
M335 VSS WL<59> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-7505 $D=0
M336 VSS WL<58> 346 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-5970 $D=0
M337 VSS WL<57> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-4435 $D=0
M338 VSS WL<56> 347 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-2900 $D=0
M339 VSS WL<55> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-1365 $D=0
M340 VSS WL<54> 348 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=170 $D=0
M341 VSS WL<53> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=1705 $D=0
M342 VSS WL<52> 349 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=3240 $D=0
M343 VSS WL<51> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=4775 $D=0
M344 VSS WL<50> 350 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=6310 $D=0
M345 VSS WL<49> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=7845 $D=0
M346 VSS WL<48> 351 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=9380 $D=0
M347 VSS WL<47> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=11335 $D=0
M348 VSS WL<46> 352 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=12870 $D=0
M349 VSS WL<45> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=14405 $D=0
M350 VSS WL<44> 353 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=15940 $D=0
M351 VSS WL<43> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=17475 $D=0
M352 VSS WL<42> 354 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=19010 $D=0
M353 VSS WL<41> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=20545 $D=0
M354 VSS WL<40> 355 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=22080 $D=0
M355 VSS WL<39> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=23615 $D=0
M356 VSS WL<38> 356 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=25150 $D=0
M357 VSS WL<37> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=26685 $D=0
M358 VSS WL<36> 357 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=28220 $D=0
M359 VSS WL<35> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=29755 $D=0
M360 VSS WL<34> 358 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=31290 $D=0
M361 VSS WL<33> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=32825 $D=0
M362 VSS WL<32> 359 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=34360 $D=0
M363 VSS WL<31> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=36315 $D=0
M364 VSS WL<30> 360 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=37850 $D=0
M365 VSS WL<29> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=39385 $D=0
M366 VSS WL<28> 361 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=40920 $D=0
M367 VSS WL<27> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=42455 $D=0
M368 VSS WL<26> 362 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=43990 $D=0
M369 VSS WL<25> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=45525 $D=0
M370 VSS WL<24> 363 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=47060 $D=0
M371 VSS WL<23> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=48595 $D=0
M372 VSS WL<22> 364 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=50130 $D=0
M373 VSS WL<21> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=51665 $D=0
M374 VSS WL<20> 365 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=53200 $D=0
M375 VSS WL<19> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=54735 $D=0
M376 VSS WL<18> 366 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=56270 $D=0
M377 VSS WL<17> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=57805 $D=0
M378 VSS WL<16> 367 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=59340 $D=0
M379 VSS WL<15> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=61295 $D=0
M380 VSS WL<14> 368 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=62830 $D=0
M381 VSS WL<13> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=64365 $D=0
M382 VSS WL<12> 369 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=65900 $D=0
M383 VSS WL<11> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=67435 $D=0
M384 VSS WL<10> 370 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=68970 $D=0
M385 VSS WL<9> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=70505 $D=0
M386 VSS WL<8> 371 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=72040 $D=0
M387 VSS WL<7> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=73575 $D=0
M388 VSS WL<6> 372 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=75110 $D=0
M389 VSS WL<5> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=76645 $D=0
M390 VSS WL<4> 373 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=78180 $D=0
M391 VSS WL<3> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=79715 $D=0
M392 VSS WL<2> 374 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=81250 $D=0
M393 VSS WL<1> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=82785 $D=0
M394 VSS WL<0> 375 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=84320 $D=0
M395 41 YOUT<3> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-25164 $Y=-35060 $D=0
M396 42 YOUT<2> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-25164 $Y=-25360 $D=0
M397 155 41 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-24979 $Y=-37026 $D=0
M398 BL<2> 42 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-24979 $Y=-27326 $D=0
M399 376 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-13645 $D=0
M400 BL<3> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-12110 $D=0
M401 377 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-10575 $D=0
M402 BL<3> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-9040 $D=0
M403 378 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-7505 $D=0
M404 BL<3> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-5970 $D=0
M405 379 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-4435 $D=0
M406 BL<3> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-2900 $D=0
M407 380 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-1365 $D=0
M408 BL<3> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=170 $D=0
M409 381 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=1705 $D=0
M410 BL<3> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=3240 $D=0
M411 382 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=4775 $D=0
M412 BL<3> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=6310 $D=0
M413 383 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=7845 $D=0
M414 BL<3> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=9380 $D=0
M415 384 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=11335 $D=0
M416 BL<3> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=12870 $D=0
M417 385 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=14405 $D=0
M418 BL<3> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=15940 $D=0
M419 386 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=17475 $D=0
M420 BL<3> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=19010 $D=0
M421 387 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=20545 $D=0
M422 BL<3> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=22080 $D=0
M423 388 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=23615 $D=0
M424 BL<3> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=25150 $D=0
M425 389 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=26685 $D=0
M426 BL<3> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=28220 $D=0
M427 390 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=29755 $D=0
M428 BL<3> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=31290 $D=0
M429 391 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=32825 $D=0
M430 BL<3> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=34360 $D=0
M431 392 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=36315 $D=0
M432 BL<3> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=37850 $D=0
M433 393 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=39385 $D=0
M434 BL<3> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=40920 $D=0
M435 394 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=42455 $D=0
M436 BL<3> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=43990 $D=0
M437 395 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=45525 $D=0
M438 BL<3> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=47060 $D=0
M439 396 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=48595 $D=0
M440 BL<3> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=50130 $D=0
M441 397 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=51665 $D=0
M442 BL<3> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=53200 $D=0
M443 398 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=54735 $D=0
M444 BL<3> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=56270 $D=0
M445 399 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=57805 $D=0
M446 BL<3> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=59340 $D=0
M447 400 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=61295 $D=0
M448 BL<3> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=62830 $D=0
M449 401 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=64365 $D=0
M450 BL<3> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=65900 $D=0
M451 402 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=67435 $D=0
M452 BL<3> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=68970 $D=0
M453 403 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=70505 $D=0
M454 BL<3> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=72040 $D=0
M455 404 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=73575 $D=0
M456 BL<3> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=75110 $D=0
M457 405 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=76645 $D=0
M458 BL<3> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=78180 $D=0
M459 406 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=79715 $D=0
M460 BL<3> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=81250 $D=0
M461 407 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=82785 $D=0
M462 BL<3> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=84320 $D=0
M463 VSS WL<63> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-13645 $D=0
M464 VSS WL<62> 408 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-12110 $D=0
M465 VSS WL<61> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-10575 $D=0
M466 VSS WL<60> 409 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-9040 $D=0
M467 VSS WL<59> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-7505 $D=0
M468 VSS WL<58> 410 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-5970 $D=0
M469 VSS WL<57> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-4435 $D=0
M470 VSS WL<56> 411 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-2900 $D=0
M471 VSS WL<55> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-1365 $D=0
M472 VSS WL<54> 412 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=170 $D=0
M473 VSS WL<53> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=1705 $D=0
M474 VSS WL<52> 413 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=3240 $D=0
M475 VSS WL<51> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=4775 $D=0
M476 VSS WL<50> 414 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=6310 $D=0
M477 VSS WL<49> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=7845 $D=0
M478 VSS WL<48> 415 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=9380 $D=0
M479 VSS WL<47> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=11335 $D=0
M480 VSS WL<46> 416 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=12870 $D=0
M481 VSS WL<45> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=14405 $D=0
M482 VSS WL<44> 417 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=15940 $D=0
M483 VSS WL<43> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=17475 $D=0
M484 VSS WL<42> 418 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=19010 $D=0
M485 VSS WL<41> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=20545 $D=0
M486 VSS WL<40> 419 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=22080 $D=0
M487 VSS WL<39> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=23615 $D=0
M488 VSS WL<38> 420 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=25150 $D=0
M489 VSS WL<37> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=26685 $D=0
M490 VSS WL<36> 421 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=28220 $D=0
M491 VSS WL<35> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=29755 $D=0
M492 VSS WL<34> 422 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=31290 $D=0
M493 VSS WL<33> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=32825 $D=0
M494 VSS WL<32> 423 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=34360 $D=0
M495 VSS WL<31> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=36315 $D=0
M496 VSS WL<30> 424 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=37850 $D=0
M497 VSS WL<29> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=39385 $D=0
M498 VSS WL<28> 425 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=40920 $D=0
M499 VSS WL<27> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=42455 $D=0
M500 VSS WL<26> 426 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=43990 $D=0
M501 VSS WL<25> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=45525 $D=0
M502 VSS WL<24> 427 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=47060 $D=0
M503 VSS WL<23> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=48595 $D=0
M504 VSS WL<22> 428 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=50130 $D=0
M505 VSS WL<21> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=51665 $D=0
M506 VSS WL<20> 429 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=53200 $D=0
M507 VSS WL<19> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=54735 $D=0
M508 VSS WL<18> 430 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=56270 $D=0
M509 VSS WL<17> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=57805 $D=0
M510 VSS WL<16> 431 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=59340 $D=0
M511 VSS WL<15> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=61295 $D=0
M512 VSS WL<14> 432 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=62830 $D=0
M513 VSS WL<13> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=64365 $D=0
M514 VSS WL<12> 433 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=65900 $D=0
M515 VSS WL<11> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=67435 $D=0
M516 VSS WL<10> 434 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=68970 $D=0
M517 VSS WL<9> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=70505 $D=0
M518 VSS WL<8> 435 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=72040 $D=0
M519 VSS WL<7> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=73575 $D=0
M520 VSS WL<6> 436 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=75110 $D=0
M521 VSS WL<5> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=76645 $D=0
M522 VSS WL<4> 437 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=78180 $D=0
M523 VSS WL<3> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=79715 $D=0
M524 VSS WL<2> 438 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=81250 $D=0
M525 VSS WL<1> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=82785 $D=0
M526 VSS WL<0> 439 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=84320 $D=0
M527 46 YOUT<5> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-23014 $Y=-35060 $D=0
M528 47 YOUT<4> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-23014 $Y=-25360 $D=0
M529 156 46 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-22829 $Y=-37026 $D=0
M530 BL<4> 47 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-22829 $Y=-27326 $D=0
M531 440 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-13645 $D=0
M532 BL<5> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-12110 $D=0
M533 441 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-10575 $D=0
M534 BL<5> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-9040 $D=0
M535 442 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-7505 $D=0
M536 BL<5> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-5970 $D=0
M537 443 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-4435 $D=0
M538 BL<5> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-2900 $D=0
M539 444 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-1365 $D=0
M540 BL<5> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=170 $D=0
M541 445 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=1705 $D=0
M542 BL<5> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=3240 $D=0
M543 446 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=4775 $D=0
M544 BL<5> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=6310 $D=0
M545 447 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=7845 $D=0
M546 BL<5> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=9380 $D=0
M547 448 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=11335 $D=0
M548 BL<5> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=12870 $D=0
M549 449 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=14405 $D=0
M550 BL<5> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=15940 $D=0
M551 450 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=17475 $D=0
M552 BL<5> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=19010 $D=0
M553 451 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=20545 $D=0
M554 BL<5> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=22080 $D=0
M555 452 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=23615 $D=0
M556 BL<5> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=25150 $D=0
M557 453 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=26685 $D=0
M558 BL<5> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=28220 $D=0
M559 454 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=29755 $D=0
M560 BL<5> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=31290 $D=0
M561 455 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=32825 $D=0
M562 BL<5> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=34360 $D=0
M563 456 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=36315 $D=0
M564 BL<5> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=37850 $D=0
M565 457 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=39385 $D=0
M566 BL<5> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=40920 $D=0
M567 458 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=42455 $D=0
M568 BL<5> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=43990 $D=0
M569 459 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=45525 $D=0
M570 BL<5> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=47060 $D=0
M571 460 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=48595 $D=0
M572 BL<5> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=50130 $D=0
M573 461 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=51665 $D=0
M574 BL<5> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=53200 $D=0
M575 462 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=54735 $D=0
M576 BL<5> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=56270 $D=0
M577 463 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=57805 $D=0
M578 BL<5> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=59340 $D=0
M579 464 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=61295 $D=0
M580 BL<5> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=62830 $D=0
M581 465 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=64365 $D=0
M582 BL<5> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=65900 $D=0
M583 466 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=67435 $D=0
M584 BL<5> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=68970 $D=0
M585 467 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=70505 $D=0
M586 BL<5> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=72040 $D=0
M587 468 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=73575 $D=0
M588 BL<5> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=75110 $D=0
M589 469 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=76645 $D=0
M590 BL<5> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=78180 $D=0
M591 470 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=79715 $D=0
M592 BL<5> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=81250 $D=0
M593 471 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=82785 $D=0
M594 BL<5> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=84320 $D=0
M595 VSS WL<63> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-13645 $D=0
M596 VSS WL<62> 472 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-12110 $D=0
M597 VSS WL<61> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-10575 $D=0
M598 VSS WL<60> 473 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-9040 $D=0
M599 VSS WL<59> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-7505 $D=0
M600 VSS WL<58> 474 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-5970 $D=0
M601 VSS WL<57> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-4435 $D=0
M602 VSS WL<56> 475 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-2900 $D=0
M603 VSS WL<55> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-1365 $D=0
M604 VSS WL<54> 476 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=170 $D=0
M605 VSS WL<53> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=1705 $D=0
M606 VSS WL<52> 477 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=3240 $D=0
M607 VSS WL<51> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=4775 $D=0
M608 VSS WL<50> 478 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=6310 $D=0
M609 VSS WL<49> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=7845 $D=0
M610 VSS WL<48> 479 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=9380 $D=0
M611 VSS WL<47> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=11335 $D=0
M612 VSS WL<46> 480 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=12870 $D=0
M613 VSS WL<45> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=14405 $D=0
M614 VSS WL<44> 481 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=15940 $D=0
M615 VSS WL<43> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=17475 $D=0
M616 VSS WL<42> 482 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=19010 $D=0
M617 VSS WL<41> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=20545 $D=0
M618 VSS WL<40> 483 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=22080 $D=0
M619 VSS WL<39> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=23615 $D=0
M620 VSS WL<38> 484 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=25150 $D=0
M621 VSS WL<37> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=26685 $D=0
M622 VSS WL<36> 485 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=28220 $D=0
M623 VSS WL<35> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=29755 $D=0
M624 VSS WL<34> 486 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=31290 $D=0
M625 VSS WL<33> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=32825 $D=0
M626 VSS WL<32> 487 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=34360 $D=0
M627 VSS WL<31> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=36315 $D=0
M628 VSS WL<30> 488 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=37850 $D=0
M629 VSS WL<29> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=39385 $D=0
M630 VSS WL<28> 489 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=40920 $D=0
M631 VSS WL<27> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=42455 $D=0
M632 VSS WL<26> 490 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=43990 $D=0
M633 VSS WL<25> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=45525 $D=0
M634 VSS WL<24> 491 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=47060 $D=0
M635 VSS WL<23> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=48595 $D=0
M636 VSS WL<22> 492 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=50130 $D=0
M637 VSS WL<21> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=51665 $D=0
M638 VSS WL<20> 493 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=53200 $D=0
M639 VSS WL<19> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=54735 $D=0
M640 VSS WL<18> 494 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=56270 $D=0
M641 VSS WL<17> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=57805 $D=0
M642 VSS WL<16> 495 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=59340 $D=0
M643 VSS WL<15> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=61295 $D=0
M644 VSS WL<14> 496 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=62830 $D=0
M645 VSS WL<13> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=64365 $D=0
M646 VSS WL<12> 497 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=65900 $D=0
M647 VSS WL<11> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=67435 $D=0
M648 VSS WL<10> 498 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=68970 $D=0
M649 VSS WL<9> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=70505 $D=0
M650 VSS WL<8> 499 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=72040 $D=0
M651 VSS WL<7> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=73575 $D=0
M652 VSS WL<6> 500 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=75110 $D=0
M653 VSS WL<5> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=76645 $D=0
M654 VSS WL<4> 501 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=78180 $D=0
M655 VSS WL<3> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=79715 $D=0
M656 VSS WL<2> 502 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=81250 $D=0
M657 VSS WL<1> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=82785 $D=0
M658 VSS WL<0> 503 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=84320 $D=0
M659 51 YOUT<7> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20864 $Y=-35060 $D=0
M660 52 YOUT<6> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20864 $Y=-25360 $D=0
M661 157 51 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20679 $Y=-37026 $D=0
M662 BL<6> 52 DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20679 $Y=-27326 $D=0
M663 504 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-13645 $D=0
M664 BL<7> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-12110 $D=0
M665 505 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-10575 $D=0
M666 BL<7> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-9040 $D=0
M667 506 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-7505 $D=0
M668 BL<7> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-5970 $D=0
M669 507 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-4435 $D=0
M670 BL<7> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-2900 $D=0
M671 508 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-1365 $D=0
M672 BL<7> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=170 $D=0
M673 509 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=1705 $D=0
M674 BL<7> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=3240 $D=0
M675 510 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=4775 $D=0
M676 BL<7> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=6310 $D=0
M677 511 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=7845 $D=0
M678 BL<7> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=9380 $D=0
M679 512 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=11335 $D=0
M680 BL<7> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=12870 $D=0
M681 513 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=14405 $D=0
M682 BL<7> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=15940 $D=0
M683 514 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=17475 $D=0
M684 BL<7> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=19010 $D=0
M685 515 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=20545 $D=0
M686 BL<7> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=22080 $D=0
M687 516 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=23615 $D=0
M688 BL<7> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=25150 $D=0
M689 517 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=26685 $D=0
M690 BL<7> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=28220 $D=0
M691 518 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=29755 $D=0
M692 BL<7> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=31290 $D=0
M693 519 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=32825 $D=0
M694 BL<7> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=34360 $D=0
M695 520 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=36315 $D=0
M696 BL<7> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=37850 $D=0
M697 521 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=39385 $D=0
M698 BL<7> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=40920 $D=0
M699 522 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=42455 $D=0
M700 BL<7> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=43990 $D=0
M701 523 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=45525 $D=0
M702 BL<7> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=47060 $D=0
M703 524 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=48595 $D=0
M704 BL<7> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=50130 $D=0
M705 525 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=51665 $D=0
M706 BL<7> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=53200 $D=0
M707 526 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=54735 $D=0
M708 BL<7> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=56270 $D=0
M709 527 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=57805 $D=0
M710 BL<7> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=59340 $D=0
M711 528 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=61295 $D=0
M712 BL<7> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=62830 $D=0
M713 529 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=64365 $D=0
M714 BL<7> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=65900 $D=0
M715 530 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=67435 $D=0
M716 BL<7> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=68970 $D=0
M717 531 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=70505 $D=0
M718 BL<7> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=72040 $D=0
M719 532 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=73575 $D=0
M720 BL<7> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=75110 $D=0
M721 533 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=76645 $D=0
M722 BL<7> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=78180 $D=0
M723 534 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=79715 $D=0
M724 BL<7> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=81250 $D=0
M725 535 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=82785 $D=0
M726 BL<7> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=84320 $D=0
M727 VSS WL<63> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-13645 $D=0
M728 VSS WL<62> 536 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-12110 $D=0
M729 VSS WL<61> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-10575 $D=0
M730 VSS WL<60> 537 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-9040 $D=0
M731 VSS WL<59> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-7505 $D=0
M732 VSS WL<58> 538 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-5970 $D=0
M733 VSS WL<57> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-4435 $D=0
M734 VSS WL<56> 539 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-2900 $D=0
M735 VSS WL<55> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-1365 $D=0
M736 VSS WL<54> 540 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=170 $D=0
M737 VSS WL<53> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=1705 $D=0
M738 VSS WL<52> 541 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=3240 $D=0
M739 VSS WL<51> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=4775 $D=0
M740 VSS WL<50> 542 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=6310 $D=0
M741 VSS WL<49> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=7845 $D=0
M742 VSS WL<48> 543 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=9380 $D=0
M743 VSS WL<47> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=11335 $D=0
M744 VSS WL<46> 544 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=12870 $D=0
M745 VSS WL<45> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=14405 $D=0
M746 VSS WL<44> 545 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=15940 $D=0
M747 VSS WL<43> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=17475 $D=0
M748 VSS WL<42> 546 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=19010 $D=0
M749 VSS WL<41> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=20545 $D=0
M750 VSS WL<40> 547 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=22080 $D=0
M751 VSS WL<39> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=23615 $D=0
M752 VSS WL<38> 548 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=25150 $D=0
M753 VSS WL<37> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=26685 $D=0
M754 VSS WL<36> 549 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=28220 $D=0
M755 VSS WL<35> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=29755 $D=0
M756 VSS WL<34> 550 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=31290 $D=0
M757 VSS WL<33> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=32825 $D=0
M758 VSS WL<32> 551 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=34360 $D=0
M759 VSS WL<31> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=36315 $D=0
M760 VSS WL<30> 552 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=37850 $D=0
M761 VSS WL<29> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=39385 $D=0
M762 VSS WL<28> 553 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=40920 $D=0
M763 VSS WL<27> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=42455 $D=0
M764 VSS WL<26> 554 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=43990 $D=0
M765 VSS WL<25> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=45525 $D=0
M766 VSS WL<24> 555 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=47060 $D=0
M767 VSS WL<23> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=48595 $D=0
M768 VSS WL<22> 556 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=50130 $D=0
M769 VSS WL<21> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=51665 $D=0
M770 VSS WL<20> 557 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=53200 $D=0
M771 VSS WL<19> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=54735 $D=0
M772 VSS WL<18> 558 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=56270 $D=0
M773 VSS WL<17> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=57805 $D=0
M774 VSS WL<16> 559 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=59340 $D=0
M775 VSS WL<15> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=61295 $D=0
M776 VSS WL<14> 560 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=62830 $D=0
M777 VSS WL<13> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=64365 $D=0
M778 VSS WL<12> 561 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=65900 $D=0
M779 VSS WL<11> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=67435 $D=0
M780 VSS WL<10> 562 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=68970 $D=0
M781 VSS WL<9> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=70505 $D=0
M782 VSS WL<8> 563 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=72040 $D=0
M783 VSS WL<7> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=73575 $D=0
M784 VSS WL<6> 564 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=75110 $D=0
M785 VSS WL<5> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=76645 $D=0
M786 VSS WL<4> 565 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=78180 $D=0
M787 VSS WL<3> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=79715 $D=0
M788 VSS WL<2> 566 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=81250 $D=0
M789 VSS WL<1> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=82785 $D=0
M790 VSS WL<0> 567 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=84320 $D=0
M791 56 YOUT<1> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18714 $Y=-35060 $D=0
M792 57 YOUT<0> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18714 $Y=-25360 $D=0
M793 159 56 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18529 $Y=-37026 $D=0
M794 BL<8> 57 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18529 $Y=-27326 $D=0
M795 568 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-13645 $D=0
M796 BL<9> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-12110 $D=0
M797 569 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-10575 $D=0
M798 BL<9> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-9040 $D=0
M799 570 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-7505 $D=0
M800 BL<9> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-5970 $D=0
M801 571 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-4435 $D=0
M802 BL<9> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-2900 $D=0
M803 572 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-1365 $D=0
M804 BL<9> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=170 $D=0
M805 573 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=1705 $D=0
M806 BL<9> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=3240 $D=0
M807 574 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=4775 $D=0
M808 BL<9> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=6310 $D=0
M809 575 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=7845 $D=0
M810 BL<9> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=9380 $D=0
M811 576 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=11335 $D=0
M812 BL<9> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=12870 $D=0
M813 577 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=14405 $D=0
M814 BL<9> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=15940 $D=0
M815 578 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=17475 $D=0
M816 BL<9> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=19010 $D=0
M817 579 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=20545 $D=0
M818 BL<9> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=22080 $D=0
M819 580 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=23615 $D=0
M820 BL<9> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=25150 $D=0
M821 581 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=26685 $D=0
M822 BL<9> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=28220 $D=0
M823 582 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=29755 $D=0
M824 BL<9> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=31290 $D=0
M825 583 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=32825 $D=0
M826 BL<9> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=34360 $D=0
M827 584 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=36315 $D=0
M828 BL<9> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=37850 $D=0
M829 585 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=39385 $D=0
M830 BL<9> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=40920 $D=0
M831 586 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=42455 $D=0
M832 BL<9> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=43990 $D=0
M833 587 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=45525 $D=0
M834 BL<9> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=47060 $D=0
M835 588 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=48595 $D=0
M836 BL<9> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=50130 $D=0
M837 589 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=51665 $D=0
M838 BL<9> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=53200 $D=0
M839 590 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=54735 $D=0
M840 BL<9> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=56270 $D=0
M841 591 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=57805 $D=0
M842 BL<9> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=59340 $D=0
M843 592 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=61295 $D=0
M844 BL<9> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=62830 $D=0
M845 593 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=64365 $D=0
M846 BL<9> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=65900 $D=0
M847 594 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=67435 $D=0
M848 BL<9> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=68970 $D=0
M849 595 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=70505 $D=0
M850 BL<9> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=72040 $D=0
M851 596 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=73575 $D=0
M852 BL<9> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=75110 $D=0
M853 597 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=76645 $D=0
M854 BL<9> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=78180 $D=0
M855 598 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=79715 $D=0
M856 BL<9> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=81250 $D=0
M857 599 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=82785 $D=0
M858 BL<9> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=84320 $D=0
M859 VSS WL<63> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-13645 $D=0
M860 VSS WL<62> 600 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-12110 $D=0
M861 VSS WL<61> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-10575 $D=0
M862 VSS WL<60> 601 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-9040 $D=0
M863 VSS WL<59> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-7505 $D=0
M864 VSS WL<58> 602 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-5970 $D=0
M865 VSS WL<57> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-4435 $D=0
M866 VSS WL<56> 603 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-2900 $D=0
M867 VSS WL<55> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-1365 $D=0
M868 VSS WL<54> 604 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=170 $D=0
M869 VSS WL<53> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=1705 $D=0
M870 VSS WL<52> 605 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=3240 $D=0
M871 VSS WL<51> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=4775 $D=0
M872 VSS WL<50> 606 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=6310 $D=0
M873 VSS WL<49> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=7845 $D=0
M874 VSS WL<48> 607 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=9380 $D=0
M875 VSS WL<47> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=11335 $D=0
M876 VSS WL<46> 608 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=12870 $D=0
M877 VSS WL<45> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=14405 $D=0
M878 VSS WL<44> 609 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=15940 $D=0
M879 VSS WL<43> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=17475 $D=0
M880 VSS WL<42> 610 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=19010 $D=0
M881 VSS WL<41> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=20545 $D=0
M882 VSS WL<40> 611 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=22080 $D=0
M883 VSS WL<39> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=23615 $D=0
M884 VSS WL<38> 612 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=25150 $D=0
M885 VSS WL<37> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=26685 $D=0
M886 VSS WL<36> 613 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=28220 $D=0
M887 VSS WL<35> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=29755 $D=0
M888 VSS WL<34> 614 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=31290 $D=0
M889 VSS WL<33> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=32825 $D=0
M890 VSS WL<32> 615 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=34360 $D=0
M891 VSS WL<31> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=36315 $D=0
M892 VSS WL<30> 616 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=37850 $D=0
M893 VSS WL<29> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=39385 $D=0
M894 VSS WL<28> 617 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=40920 $D=0
M895 VSS WL<27> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=42455 $D=0
M896 VSS WL<26> 618 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=43990 $D=0
M897 VSS WL<25> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=45525 $D=0
M898 VSS WL<24> 619 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=47060 $D=0
M899 VSS WL<23> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=48595 $D=0
M900 VSS WL<22> 620 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=50130 $D=0
M901 VSS WL<21> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=51665 $D=0
M902 VSS WL<20> 621 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=53200 $D=0
M903 VSS WL<19> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=54735 $D=0
M904 VSS WL<18> 622 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=56270 $D=0
M905 VSS WL<17> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=57805 $D=0
M906 VSS WL<16> 623 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=59340 $D=0
M907 VSS WL<15> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=61295 $D=0
M908 VSS WL<14> 624 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=62830 $D=0
M909 VSS WL<13> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=64365 $D=0
M910 VSS WL<12> 625 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=65900 $D=0
M911 VSS WL<11> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=67435 $D=0
M912 VSS WL<10> 626 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=68970 $D=0
M913 VSS WL<9> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=70505 $D=0
M914 VSS WL<8> 627 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=72040 $D=0
M915 VSS WL<7> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=73575 $D=0
M916 VSS WL<6> 628 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=75110 $D=0
M917 VSS WL<5> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=76645 $D=0
M918 VSS WL<4> 629 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=78180 $D=0
M919 VSS WL<3> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=79715 $D=0
M920 VSS WL<2> 630 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=81250 $D=0
M921 VSS WL<1> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=82785 $D=0
M922 VSS WL<0> 631 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=84320 $D=0
M923 61 YOUT<3> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16564 $Y=-35060 $D=0
M924 62 YOUT<2> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16564 $Y=-25360 $D=0
M925 160 61 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16379 $Y=-37026 $D=0
M926 BL<10> 62 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16379 $Y=-27326 $D=0
M927 632 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-13645 $D=0
M928 BL<11> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-12110 $D=0
M929 633 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-10575 $D=0
M930 BL<11> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-9040 $D=0
M931 634 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-7505 $D=0
M932 BL<11> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-5970 $D=0
M933 635 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-4435 $D=0
M934 BL<11> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-2900 $D=0
M935 636 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-1365 $D=0
M936 BL<11> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=170 $D=0
M937 637 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=1705 $D=0
M938 BL<11> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=3240 $D=0
M939 638 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=4775 $D=0
M940 BL<11> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=6310 $D=0
M941 639 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=7845 $D=0
M942 BL<11> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=9380 $D=0
M943 640 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=11335 $D=0
M944 BL<11> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=12870 $D=0
M945 641 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=14405 $D=0
M946 BL<11> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=15940 $D=0
M947 642 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=17475 $D=0
M948 BL<11> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=19010 $D=0
M949 643 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=20545 $D=0
M950 BL<11> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=22080 $D=0
M951 644 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=23615 $D=0
M952 BL<11> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=25150 $D=0
M953 645 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=26685 $D=0
M954 BL<11> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=28220 $D=0
M955 646 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=29755 $D=0
M956 BL<11> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=31290 $D=0
M957 647 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=32825 $D=0
M958 BL<11> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=34360 $D=0
M959 648 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=36315 $D=0
M960 BL<11> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=37850 $D=0
M961 649 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=39385 $D=0
M962 BL<11> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=40920 $D=0
M963 650 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=42455 $D=0
M964 BL<11> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=43990 $D=0
M965 651 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=45525 $D=0
M966 BL<11> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=47060 $D=0
M967 652 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=48595 $D=0
M968 BL<11> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=50130 $D=0
M969 653 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=51665 $D=0
M970 BL<11> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=53200 $D=0
M971 654 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=54735 $D=0
M972 BL<11> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=56270 $D=0
M973 655 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=57805 $D=0
M974 BL<11> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=59340 $D=0
M975 656 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=61295 $D=0
M976 BL<11> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=62830 $D=0
M977 657 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=64365 $D=0
M978 BL<11> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=65900 $D=0
M979 658 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=67435 $D=0
M980 BL<11> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=68970 $D=0
M981 659 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=70505 $D=0
M982 BL<11> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=72040 $D=0
M983 660 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=73575 $D=0
M984 BL<11> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=75110 $D=0
M985 661 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=76645 $D=0
M986 BL<11> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=78180 $D=0
M987 662 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=79715 $D=0
M988 BL<11> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=81250 $D=0
M989 663 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=82785 $D=0
M990 BL<11> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=84320 $D=0
M991 VSS WL<63> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-13645 $D=0
M992 VSS WL<62> 664 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-12110 $D=0
M993 VSS WL<61> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-10575 $D=0
M994 VSS WL<60> 665 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-9040 $D=0
M995 VSS WL<59> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-7505 $D=0
M996 VSS WL<58> 666 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-5970 $D=0
M997 VSS WL<57> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-4435 $D=0
M998 VSS WL<56> 667 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-2900 $D=0
M999 VSS WL<55> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-1365 $D=0
M1000 VSS WL<54> 668 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=170 $D=0
M1001 VSS WL<53> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=1705 $D=0
M1002 VSS WL<52> 669 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=3240 $D=0
M1003 VSS WL<51> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=4775 $D=0
M1004 VSS WL<50> 670 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=6310 $D=0
M1005 VSS WL<49> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=7845 $D=0
M1006 VSS WL<48> 671 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=9380 $D=0
M1007 VSS WL<47> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=11335 $D=0
M1008 VSS WL<46> 672 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=12870 $D=0
M1009 VSS WL<45> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=14405 $D=0
M1010 VSS WL<44> 673 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=15940 $D=0
M1011 VSS WL<43> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=17475 $D=0
M1012 VSS WL<42> 674 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=19010 $D=0
M1013 VSS WL<41> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=20545 $D=0
M1014 VSS WL<40> 675 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=22080 $D=0
M1015 VSS WL<39> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=23615 $D=0
M1016 VSS WL<38> 676 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=25150 $D=0
M1017 VSS WL<37> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=26685 $D=0
M1018 VSS WL<36> 677 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=28220 $D=0
M1019 VSS WL<35> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=29755 $D=0
M1020 VSS WL<34> 678 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=31290 $D=0
M1021 VSS WL<33> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=32825 $D=0
M1022 VSS WL<32> 679 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=34360 $D=0
M1023 VSS WL<31> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=36315 $D=0
M1024 VSS WL<30> 680 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=37850 $D=0
M1025 VSS WL<29> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=39385 $D=0
M1026 VSS WL<28> 681 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=40920 $D=0
M1027 VSS WL<27> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=42455 $D=0
M1028 VSS WL<26> 682 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=43990 $D=0
M1029 VSS WL<25> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=45525 $D=0
M1030 VSS WL<24> 683 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=47060 $D=0
M1031 VSS WL<23> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=48595 $D=0
M1032 VSS WL<22> 684 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=50130 $D=0
M1033 VSS WL<21> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=51665 $D=0
M1034 VSS WL<20> 685 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=53200 $D=0
M1035 VSS WL<19> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=54735 $D=0
M1036 VSS WL<18> 686 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=56270 $D=0
M1037 VSS WL<17> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=57805 $D=0
M1038 VSS WL<16> 687 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=59340 $D=0
M1039 VSS WL<15> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=61295 $D=0
M1040 VSS WL<14> 688 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=62830 $D=0
M1041 VSS WL<13> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=64365 $D=0
M1042 VSS WL<12> 689 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=65900 $D=0
M1043 VSS WL<11> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=67435 $D=0
M1044 VSS WL<10> 690 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=68970 $D=0
M1045 VSS WL<9> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=70505 $D=0
M1046 VSS WL<8> 691 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=72040 $D=0
M1047 VSS WL<7> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=73575 $D=0
M1048 VSS WL<6> 692 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=75110 $D=0
M1049 VSS WL<5> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=76645 $D=0
M1050 VSS WL<4> 693 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=78180 $D=0
M1051 VSS WL<3> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=79715 $D=0
M1052 VSS WL<2> 694 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=81250 $D=0
M1053 VSS WL<1> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=82785 $D=0
M1054 VSS WL<0> 695 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=84320 $D=0
M1055 66 YOUT<5> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14414 $Y=-35060 $D=0
M1056 67 YOUT<4> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14414 $Y=-25360 $D=0
M1057 161 66 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14229 $Y=-37026 $D=0
M1058 BL<12> 67 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14229 $Y=-27326 $D=0
M1059 696 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-13645 $D=0
M1060 BL<13> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-12110 $D=0
M1061 697 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-10575 $D=0
M1062 BL<13> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-9040 $D=0
M1063 698 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-7505 $D=0
M1064 BL<13> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-5970 $D=0
M1065 699 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-4435 $D=0
M1066 BL<13> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-2900 $D=0
M1067 700 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-1365 $D=0
M1068 BL<13> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=170 $D=0
M1069 701 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=1705 $D=0
M1070 BL<13> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=3240 $D=0
M1071 702 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=4775 $D=0
M1072 BL<13> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=6310 $D=0
M1073 703 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=7845 $D=0
M1074 BL<13> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=9380 $D=0
M1075 704 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=11335 $D=0
M1076 BL<13> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=12870 $D=0
M1077 705 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=14405 $D=0
M1078 BL<13> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=15940 $D=0
M1079 706 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=17475 $D=0
M1080 BL<13> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=19010 $D=0
M1081 707 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=20545 $D=0
M1082 BL<13> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=22080 $D=0
M1083 708 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=23615 $D=0
M1084 BL<13> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=25150 $D=0
M1085 709 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=26685 $D=0
M1086 BL<13> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=28220 $D=0
M1087 710 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=29755 $D=0
M1088 BL<13> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=31290 $D=0
M1089 711 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=32825 $D=0
M1090 BL<13> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=34360 $D=0
M1091 712 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=36315 $D=0
M1092 BL<13> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=37850 $D=0
M1093 713 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=39385 $D=0
M1094 BL<13> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=40920 $D=0
M1095 714 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=42455 $D=0
M1096 BL<13> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=43990 $D=0
M1097 715 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=45525 $D=0
M1098 BL<13> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=47060 $D=0
M1099 716 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=48595 $D=0
M1100 BL<13> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=50130 $D=0
M1101 717 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=51665 $D=0
M1102 BL<13> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=53200 $D=0
M1103 718 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=54735 $D=0
M1104 BL<13> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=56270 $D=0
M1105 719 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=57805 $D=0
M1106 BL<13> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=59340 $D=0
M1107 720 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=61295 $D=0
M1108 BL<13> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=62830 $D=0
M1109 721 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=64365 $D=0
M1110 BL<13> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=65900 $D=0
M1111 722 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=67435 $D=0
M1112 BL<13> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=68970 $D=0
M1113 723 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=70505 $D=0
M1114 BL<13> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=72040 $D=0
M1115 724 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=73575 $D=0
M1116 BL<13> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=75110 $D=0
M1117 725 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=76645 $D=0
M1118 BL<13> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=78180 $D=0
M1119 726 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=79715 $D=0
M1120 BL<13> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=81250 $D=0
M1121 727 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=82785 $D=0
M1122 BL<13> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=84320 $D=0
M1123 VSS WL<63> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-13645 $D=0
M1124 VSS WL<62> 728 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-12110 $D=0
M1125 VSS WL<61> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-10575 $D=0
M1126 VSS WL<60> 729 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-9040 $D=0
M1127 VSS WL<59> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-7505 $D=0
M1128 VSS WL<58> 730 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-5970 $D=0
M1129 VSS WL<57> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-4435 $D=0
M1130 VSS WL<56> 731 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-2900 $D=0
M1131 VSS WL<55> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-1365 $D=0
M1132 VSS WL<54> 732 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=170 $D=0
M1133 VSS WL<53> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=1705 $D=0
M1134 VSS WL<52> 733 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=3240 $D=0
M1135 VSS WL<51> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=4775 $D=0
M1136 VSS WL<50> 734 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=6310 $D=0
M1137 VSS WL<49> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=7845 $D=0
M1138 VSS WL<48> 735 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=9380 $D=0
M1139 VSS WL<47> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=11335 $D=0
M1140 VSS WL<46> 736 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=12870 $D=0
M1141 VSS WL<45> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=14405 $D=0
M1142 VSS WL<44> 737 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=15940 $D=0
M1143 VSS WL<43> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=17475 $D=0
M1144 VSS WL<42> 738 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=19010 $D=0
M1145 VSS WL<41> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=20545 $D=0
M1146 VSS WL<40> 739 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=22080 $D=0
M1147 VSS WL<39> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=23615 $D=0
M1148 VSS WL<38> 740 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=25150 $D=0
M1149 VSS WL<37> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=26685 $D=0
M1150 VSS WL<36> 741 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=28220 $D=0
M1151 VSS WL<35> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=29755 $D=0
M1152 VSS WL<34> 742 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=31290 $D=0
M1153 VSS WL<33> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=32825 $D=0
M1154 VSS WL<32> 743 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=34360 $D=0
M1155 VSS WL<31> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=36315 $D=0
M1156 VSS WL<30> 744 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=37850 $D=0
M1157 VSS WL<29> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=39385 $D=0
M1158 VSS WL<28> 745 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=40920 $D=0
M1159 VSS WL<27> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=42455 $D=0
M1160 VSS WL<26> 746 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=43990 $D=0
M1161 VSS WL<25> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=45525 $D=0
M1162 VSS WL<24> 747 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=47060 $D=0
M1163 VSS WL<23> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=48595 $D=0
M1164 VSS WL<22> 748 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=50130 $D=0
M1165 VSS WL<21> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=51665 $D=0
M1166 VSS WL<20> 749 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=53200 $D=0
M1167 VSS WL<19> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=54735 $D=0
M1168 VSS WL<18> 750 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=56270 $D=0
M1169 VSS WL<17> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=57805 $D=0
M1170 VSS WL<16> 751 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=59340 $D=0
M1171 VSS WL<15> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=61295 $D=0
M1172 VSS WL<14> 752 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=62830 $D=0
M1173 VSS WL<13> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=64365 $D=0
M1174 VSS WL<12> 753 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=65900 $D=0
M1175 VSS WL<11> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=67435 $D=0
M1176 VSS WL<10> 754 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=68970 $D=0
M1177 VSS WL<9> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=70505 $D=0
M1178 VSS WL<8> 755 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=72040 $D=0
M1179 VSS WL<7> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=73575 $D=0
M1180 VSS WL<6> 756 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=75110 $D=0
M1181 VSS WL<5> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=76645 $D=0
M1182 VSS WL<4> 757 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=78180 $D=0
M1183 VSS WL<3> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=79715 $D=0
M1184 VSS WL<2> 758 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=81250 $D=0
M1185 VSS WL<1> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=82785 $D=0
M1186 VSS WL<0> 759 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=84320 $D=0
M1187 71 YOUT<7> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12264 $Y=-35060 $D=0
M1188 72 YOUT<6> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12264 $Y=-25360 $D=0
M1189 162 71 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12079 $Y=-37026 $D=0
M1190 BL<14> 72 DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12079 $Y=-27326 $D=0
M1191 760 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-13645 $D=0
M1192 BL<15> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-12110 $D=0
M1193 761 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-10575 $D=0
M1194 BL<15> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-9040 $D=0
M1195 762 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-7505 $D=0
M1196 BL<15> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-5970 $D=0
M1197 763 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-4435 $D=0
M1198 BL<15> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-2900 $D=0
M1199 764 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-1365 $D=0
M1200 BL<15> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=170 $D=0
M1201 765 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=1705 $D=0
M1202 BL<15> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=3240 $D=0
M1203 766 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=4775 $D=0
M1204 BL<15> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=6310 $D=0
M1205 767 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=7845 $D=0
M1206 BL<15> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=9380 $D=0
M1207 768 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=11335 $D=0
M1208 BL<15> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=12870 $D=0
M1209 769 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=14405 $D=0
M1210 BL<15> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=15940 $D=0
M1211 770 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=17475 $D=0
M1212 BL<15> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=19010 $D=0
M1213 771 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=20545 $D=0
M1214 BL<15> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=22080 $D=0
M1215 772 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=23615 $D=0
M1216 BL<15> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=25150 $D=0
M1217 773 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=26685 $D=0
M1218 BL<15> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=28220 $D=0
M1219 774 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=29755 $D=0
M1220 BL<15> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=31290 $D=0
M1221 775 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=32825 $D=0
M1222 BL<15> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=34360 $D=0
M1223 776 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=36315 $D=0
M1224 BL<15> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=37850 $D=0
M1225 777 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=39385 $D=0
M1226 BL<15> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=40920 $D=0
M1227 778 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=42455 $D=0
M1228 BL<15> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=43990 $D=0
M1229 779 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=45525 $D=0
M1230 BL<15> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=47060 $D=0
M1231 780 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=48595 $D=0
M1232 BL<15> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=50130 $D=0
M1233 781 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=51665 $D=0
M1234 BL<15> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=53200 $D=0
M1235 782 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=54735 $D=0
M1236 BL<15> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=56270 $D=0
M1237 783 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=57805 $D=0
M1238 BL<15> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=59340 $D=0
M1239 784 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=61295 $D=0
M1240 BL<15> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=62830 $D=0
M1241 785 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=64365 $D=0
M1242 BL<15> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=65900 $D=0
M1243 786 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=67435 $D=0
M1244 BL<15> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=68970 $D=0
M1245 787 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=70505 $D=0
M1246 BL<15> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=72040 $D=0
M1247 788 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=73575 $D=0
M1248 BL<15> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=75110 $D=0
M1249 789 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=76645 $D=0
M1250 BL<15> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=78180 $D=0
M1251 790 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=79715 $D=0
M1252 BL<15> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=81250 $D=0
M1253 791 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=82785 $D=0
M1254 BL<15> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=84320 $D=0
M1255 83 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=8965 $D=1
M1256 81 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=21005 $D=1
M1257 85 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=33045 $D=1
M1258 84 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=57645 $D=1
M1259 82 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=69685 $D=1
M1260 86 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=81725 $D=1
M1261 16 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-11510 $D=1
M1262 16 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-10050 $D=1
M1263 16 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-8590 $D=1
M1264 16 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-7130 $D=1
M1265 17 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-5490 $D=1
M1266 17 83 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-4030 $D=1
M1267 17 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-2570 $D=1
M1268 17 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-1110 $D=1
M1269 18 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=530 $D=1
M1270 18 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=1990 $D=1
M1271 18 81 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=3450 $D=1
M1272 18 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=4910 $D=1
M1273 19 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=6550 $D=1
M1274 19 83 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=8010 $D=1
M1275 19 81 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=9470 $D=1
M1276 19 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=10930 $D=1
M1277 20 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=12570 $D=1
M1278 20 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=14030 $D=1
M1279 20 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=15490 $D=1
M1280 20 85 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=16950 $D=1
M1281 21 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=18590 $D=1
M1282 21 83 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=20050 $D=1
M1283 21 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=21510 $D=1
M1284 21 85 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=22970 $D=1
M1285 22 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=24610 $D=1
M1286 22 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=26070 $D=1
M1287 22 81 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=27530 $D=1
M1288 22 85 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=28990 $D=1
M1289 23 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=30630 $D=1
M1290 23 83 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=32090 $D=1
M1291 23 81 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=33550 $D=1
M1292 23 85 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=35010 $D=1
M1293 24 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=37170 $D=1
M1294 24 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=38630 $D=1
M1295 24 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=40090 $D=1
M1296 24 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=41550 $D=1
M1297 25 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=43190 $D=1
M1298 25 84 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=44650 $D=1
M1299 25 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=46110 $D=1
M1300 25 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=47570 $D=1
M1301 26 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=49210 $D=1
M1302 26 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=50670 $D=1
M1303 26 82 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=52130 $D=1
M1304 26 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=53590 $D=1
M1305 27 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=55230 $D=1
M1306 27 84 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=56690 $D=1
M1307 27 82 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=58150 $D=1
M1308 27 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=59610 $D=1
M1309 28 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=61250 $D=1
M1310 28 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=62710 $D=1
M1311 28 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=64170 $D=1
M1312 28 86 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=65630 $D=1
M1313 29 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=67270 $D=1
M1314 29 84 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=68730 $D=1
M1315 29 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=70190 $D=1
M1316 29 86 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=71650 $D=1
M1317 30 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=73290 $D=1
M1318 30 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=74750 $D=1
M1319 30 82 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=76210 $D=1
M1320 30 86 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=77670 $D=1
M1321 31 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=79310 $D=1
M1322 31 84 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=80770 $D=1
M1323 31 82 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=82230 $D=1
M1324 31 86 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=83690 $D=1
M1325 WL<63> 16 216 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-13505 $D=1
M1326 WL<62> 16 217 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-11970 $D=1
M1327 WL<61> 16 218 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-10435 $D=1
M1328 WL<60> 16 219 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-8900 $D=1
M1329 WL<59> 16 220 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-7365 $D=1
M1330 WL<58> 16 221 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-5830 $D=1
M1331 WL<57> 16 222 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-4295 $D=1
M1332 WL<56> 16 223 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-2760 $D=1
M1333 WL<55> 17 224 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-1225 $D=1
M1334 WL<54> 17 225 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=310 $D=1
M1335 WL<53> 17 226 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=1845 $D=1
M1336 WL<52> 17 227 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=3380 $D=1
M1337 WL<51> 17 228 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=4915 $D=1
M1338 WL<50> 17 229 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=6450 $D=1
M1339 WL<49> 17 230 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=7985 $D=1
M1340 WL<48> 17 231 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=9520 $D=1
M1341 WL<47> 18 232 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=11475 $D=1
M1342 WL<46> 18 233 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=13010 $D=1
M1343 WL<45> 18 234 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=14545 $D=1
M1344 WL<44> 18 235 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=16080 $D=1
M1345 WL<43> 18 236 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=17615 $D=1
M1346 WL<42> 18 237 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=19150 $D=1
M1347 WL<41> 18 238 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=20685 $D=1
M1348 WL<40> 18 239 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=22220 $D=1
M1349 WL<39> 19 240 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=23755 $D=1
M1350 WL<38> 19 241 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=25290 $D=1
M1351 WL<37> 19 242 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=26825 $D=1
M1352 WL<36> 19 243 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=28360 $D=1
M1353 WL<35> 19 244 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=29895 $D=1
M1354 WL<34> 19 245 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=31430 $D=1
M1355 WL<33> 19 246 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=32965 $D=1
M1356 WL<32> 19 247 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=34500 $D=1
M1357 WL<31> 20 248 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=36455 $D=1
M1358 WL<30> 20 249 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=37990 $D=1
M1359 WL<29> 20 250 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=39525 $D=1
M1360 WL<28> 20 251 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=41060 $D=1
M1361 WL<27> 20 252 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=42595 $D=1
M1362 WL<26> 20 253 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=44130 $D=1
M1363 WL<25> 20 254 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=45665 $D=1
M1364 WL<24> 20 255 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=47200 $D=1
M1365 WL<23> 21 256 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=48735 $D=1
M1366 WL<22> 21 257 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=50270 $D=1
M1367 WL<21> 21 258 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=51805 $D=1
M1368 WL<20> 21 259 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=53340 $D=1
M1369 WL<19> 21 260 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=54875 $D=1
M1370 WL<18> 21 261 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=56410 $D=1
M1371 WL<17> 21 262 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=57945 $D=1
M1372 WL<16> 21 263 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=59480 $D=1
M1373 WL<15> 22 264 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=61435 $D=1
M1374 WL<14> 22 265 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=62970 $D=1
M1375 WL<13> 22 266 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=64505 $D=1
M1376 WL<12> 22 267 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=66040 $D=1
M1377 WL<11> 22 268 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=67575 $D=1
M1378 WL<10> 22 269 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=69110 $D=1
M1379 WL<9> 22 270 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=70645 $D=1
M1380 WL<8> 22 271 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=72180 $D=1
M1381 WL<7> 23 272 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=73715 $D=1
M1382 WL<6> 23 273 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=75250 $D=1
M1383 WL<5> 23 274 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=76785 $D=1
M1384 WL<4> 23 275 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=78320 $D=1
M1385 WL<3> 23 276 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=79855 $D=1
M1386 WL<2> 23 277 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=81390 $D=1
M1387 WL<1> 23 278 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=82925 $D=1
M1388 WL<0> 23 279 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=84460 $D=1
M1389 VDD 24 216 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-13505 $D=1
M1390 VDD 25 217 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-11970 $D=1
M1391 VDD 26 218 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-10435 $D=1
M1392 VDD 27 219 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-8900 $D=1
M1393 VDD 28 220 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-7365 $D=1
M1394 VDD 29 221 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-5830 $D=1
M1395 VDD 30 222 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-4295 $D=1
M1396 VDD 31 223 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-2760 $D=1
M1397 VDD 24 224 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-1225 $D=1
M1398 VDD 25 225 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=310 $D=1
M1399 VDD 26 226 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=1845 $D=1
M1400 VDD 27 227 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=3380 $D=1
M1401 VDD 28 228 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=4915 $D=1
M1402 VDD 29 229 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=6450 $D=1
M1403 VDD 30 230 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=7985 $D=1
M1404 VDD 31 231 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=9520 $D=1
M1405 VDD 24 232 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=11475 $D=1
M1406 VDD 25 233 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=13010 $D=1
M1407 VDD 26 234 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=14545 $D=1
M1408 VDD 27 235 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=16080 $D=1
M1409 VDD 28 236 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=17615 $D=1
M1410 VDD 29 237 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=19150 $D=1
M1411 VDD 30 238 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=20685 $D=1
M1412 VDD 31 239 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=22220 $D=1
M1413 VDD 24 240 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=23755 $D=1
M1414 VDD 25 241 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=25290 $D=1
M1415 VDD 26 242 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=26825 $D=1
M1416 VDD 27 243 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=28360 $D=1
M1417 VDD 28 244 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=29895 $D=1
M1418 VDD 29 245 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=31430 $D=1
M1419 VDD 30 246 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=32965 $D=1
M1420 VDD 31 247 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=34500 $D=1
M1421 VDD 24 248 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=36455 $D=1
M1422 VDD 25 249 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=37990 $D=1
M1423 VDD 26 250 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=39525 $D=1
M1424 VDD 27 251 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=41060 $D=1
M1425 VDD 28 252 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=42595 $D=1
M1426 VDD 29 253 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=44130 $D=1
M1427 VDD 30 254 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=45665 $D=1
M1428 VDD 31 255 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=47200 $D=1
M1429 VDD 24 256 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=48735 $D=1
M1430 VDD 25 257 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=50270 $D=1
M1431 VDD 26 258 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=51805 $D=1
M1432 VDD 27 259 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=53340 $D=1
M1433 VDD 28 260 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=54875 $D=1
M1434 VDD 29 261 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=56410 $D=1
M1435 VDD 30 262 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=57945 $D=1
M1436 VDD 31 263 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=59480 $D=1
M1437 VDD 24 264 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=61435 $D=1
M1438 VDD 25 265 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=62970 $D=1
M1439 VDD 26 266 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=64505 $D=1
M1440 VDD 27 267 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=66040 $D=1
M1441 VDD 28 268 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=67575 $D=1
M1442 VDD 29 269 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=69110 $D=1
M1443 VDD 30 270 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=70645 $D=1
M1444 VDD 31 271 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=72180 $D=1
M1445 VDD 24 272 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=73715 $D=1
M1446 VDD 25 273 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=75250 $D=1
M1447 VDD 26 274 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=76785 $D=1
M1448 VDD 27 275 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=78320 $D=1
M1449 VDD 28 276 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=79855 $D=1
M1450 VDD 29 277 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=81390 $D=1
M1451 VDD 30 278 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=82925 $D=1
M1452 VDD 31 279 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=84460 $D=1
M1453 VDD CLK BL<0> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-27660 $Y=-17045 $D=1
M1454 36 YOUT<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-33355 $D=1
M1455 DL<0> YOUT<1> 154 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-30455 $D=1
M1456 37 YOUT<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-23655 $D=1
M1457 DL<0> YOUT<0> BL<0> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-20755 $D=1
M1458 BL<1> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-26970 $Y=-17045 $D=1
M1459 VDD CLK BL<2> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-25510 $Y=-17045 $D=1
M1460 42 YOUT<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-25164 $Y=-23655 $D=1
M1461 DL<0> YOUT<2> BL<2> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-25164 $Y=-20755 $D=1
M1462 BL<3> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-24820 $Y=-17045 $D=1
M1463 VDD CLK BL<4> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-23360 $Y=-17045 $D=1
M1464 46 YOUT<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-33355 $D=1
M1465 DL<0> YOUT<5> 156 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-30455 $D=1
M1466 47 YOUT<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-23655 $D=1
M1467 DL<0> YOUT<4> BL<4> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-20755 $D=1
M1468 BL<5> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-22670 $Y=-17045 $D=1
M1469 VDD CLK BL<6> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-21210 $Y=-17045 $D=1
M1470 51 YOUT<7> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-33355 $D=1
M1471 DL<0> YOUT<7> 157 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-30455 $D=1
M1472 52 YOUT<6> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-23655 $D=1
M1473 DL<0> YOUT<6> BL<6> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-20755 $D=1
M1474 BL<7> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-20520 $Y=-17045 $D=1
M1475 VDD CLK BL<8> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-19060 $Y=-17045 $D=1
M1476 56 YOUT<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-33355 $D=1
M1477 DL<1> YOUT<1> 159 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-30455 $D=1
M1478 57 YOUT<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-23655 $D=1
M1479 DL<1> YOUT<0> BL<8> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-20755 $D=1
M1480 BL<9> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-18370 $Y=-17045 $D=1
M1481 VDD CLK BL<10> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-16910 $Y=-17045 $D=1
M1482 61 YOUT<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-33355 $D=1
M1483 DL<1> YOUT<3> 160 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-30455 $D=1
M1484 62 YOUT<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-23655 $D=1
M1485 DL<1> YOUT<2> BL<10> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-20755 $D=1
M1486 BL<11> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-16220 $Y=-17045 $D=1
M1487 VDD CLK BL<12> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-14760 $Y=-17045 $D=1
M1488 66 YOUT<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-33355 $D=1
M1489 DL<1> YOUT<5> 161 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-30455 $D=1
M1490 67 YOUT<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-23655 $D=1
M1491 DL<1> YOUT<4> BL<12> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-20755 $D=1
M1492 BL<13> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-14070 $Y=-17045 $D=1
M1493 VDD CLK BL<14> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-12610 $Y=-17045 $D=1
M1494 71 YOUT<7> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-33355 $D=1
M1495 DL<1> YOUT<7> 162 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-30455 $D=1
M1496 72 YOUT<6> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-23655 $D=1
M1497 DL<1> YOUT<6> BL<14> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-20755 $D=1
M1498 BL<15> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-11920 $Y=-17045 $D=1
X1499 Dout<0> SO<0> SAEN DL<0> VSS Vref VDD Final_SA $T=-23415 -43080 0 0 $X=-26580 $Y=-45535
X1500 Dout<1> SO<1> SAEN DL<1> VSS Vref VDD Final_SA $T=-15255 -43080 0 0 $X=-18420 $Y=-45535
X1501 CLK VSS VDD 9 inv_final $T=-68030 -26395 0 0 $X=-69190 $Y=-29660
X1502 793 VSS VDD 165 inv_final $T=-65830 -33650 0 0 $X=-66990 $Y=-36915
X1503 CLK 88 VDD VSS WL_EN final_and $T=-60940 -45770 0 0 $X=-54185 $Y=-46920
X1504 CLK 89 VDD VSS SAEN final_and $T=-48650 -45770 0 0 $X=-41895 $Y=-46920
X1505 Y_sel<0> Y_sel<1> Y_sel<2> YOUT<3> YOUT<2> YOUT<1> YOUT<0> YOUT<7> YOUT<6> YOUT<5> YOUT<4> VDD VSS Ydecoder_final $T=-62410 -36975 0 0 $X=-62790 $Y=-40160
X1506 794 VSS VDD 795 793 ICV_2 $T=-69030 -33650 0 0 $X=-70190 $Y=-36915
X1507 796 VSS VDD 797 794 ICV_3 $T=-75430 -33650 0 0 $X=-76590 $Y=-36915
X1508 798 VSS VDD 799 87 ICV_3 $T=-62670 -43335 0 0 $X=-63830 $Y=-46600
X1509 800 VSS VDD 89 88 ICV_3 $T=-62475 -50525 0 0 $X=-63635 $Y=-53790
X1510 165 VSS VDD 801 ICV_4 $T=-88270 -43335 0 0 $X=-89430 $Y=-46600
X1511 CLK VSS VDD 796 ICV_4 $T=-88230 -33650 0 0 $X=-89390 $Y=-36915
X1512 87 VSS VDD 802 ICV_4 $T=-88075 -50525 0 0 $X=-89235 $Y=-53790
X1513 801 VSS VDD 798 ICV_4 $T=-75470 -43335 0 0 $X=-76630 $Y=-46600
X1514 802 VSS VDD 800 ICV_4 $T=-75275 -50525 0 0 $X=-76435 $Y=-53790
X1515 9 CLK VSS VDD A<2> Y_sel<2> FInal_FF $T=-84440 -21020 0 0 $X=-90065 $Y=-28235
X1516 9 CLK VSS VDD A<1> Y_sel<1> FInal_FF $T=-84440 -8310 0 0 $X=-90065 $Y=-15525
X1517 9 CLK VSS VDD A<0> Y_sel<0> FInal_FF $T=-84440 4400 0 0 $X=-90065 $Y=-2815
X1518 9 CLK VSS VDD A<6> X_sel<3> FInal_FF $T=-84440 17110 0 0 $X=-90065 $Y=9895
X1519 9 CLK VSS VDD A<7> X_sel<4> FInal_FF $T=-84440 29820 0 0 $X=-90065 $Y=22605
X1520 9 CLK VSS VDD A<8> X_sel<5> FInal_FF $T=-84440 42530 0 0 $X=-90065 $Y=35315
X1521 9 CLK VSS VDD A<3> X_sel<0> FInal_FF $T=-84440 55240 0 0 $X=-90065 $Y=48025
X1522 9 CLK VSS VDD A<4> X_sel<1> FInal_FF $T=-84440 67950 0 0 $X=-90065 $Y=60735
X1523 9 CLK VSS VDD A<5> X_sel<2> FInal_FF $T=-84440 80660 0 0 $X=-90065 $Y=73445
*.CALIBRE WARNING SCONNECT SCONNECT conflict(s) detected by extraction in this cell. See extraction report for details.
** WARNING: BAD DEVICE on layer PG_SP at location (-25.164,-33.355) in cell Final_all_v1 (see extraction report).
*.CALIBRE WARNING BADDEV BAD DEVICE(s) detected by extraction in this cell. See extraction report for details.
** WARNING: BAD DEVICE on layer PG_SP at location (-25.164,-30.455) in cell Final_all_v1 (see extraction report).
.ENDS
***************************************
