************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: inverter
* View Name:     schematic
* Netlisted on:  Jan  5 12:22:19 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter IN OUT VDD VSS
*.PININFO IN:I OUT:B VDD:B VSS:B
MM10 OUT IN VSS VSS NM W=500.0n L=180.00n m=1
MM6 OUT IN VDD VDD PM W=2u L=180.00n m=1
.ENDS

