* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT pmos_small
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1
** N=5 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4
** N=5 EP=4 IP=14 FDC=1
M0 2 3 1 4 P_18 L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=1.225e-12 PD=3.48e-06 PS=3.48e-06 $X=-3180 $Y=-1840 $D=1
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4
** N=5 EP=4 IP=10 FDC=2
X0 1 2 3 4 ICV_2 $T=-1460 0 0 0 $X=-5630 $Y=-3490
X1 1 2 3 4 ICV_2 $T=0 0 0 0 $X=-4170 $Y=-3490
.ENDS
***************************************
.SUBCKT ICV_4
** N=4 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3
** N=4 EP=3 IP=12 FDC=1
M0 2 3 1 2 P_18 L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=1.225e-12 PD=3.48e-06 PS=3.48e-06 $X=-3180 $Y=160 $D=1
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3
** N=4 EP=3 IP=8 FDC=2
X0 1 2 3 ICV_5 $T=0 0 0 0 $X=-4170 $Y=-1490
X1 1 2 3 ICV_5 $T=1460 0 0 0 $X=-2710 $Y=-1490
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3
** N=4 EP=3 IP=8 FDC=4
X0 1 2 3 ICV_6 $T=0 0 0 0 $X=-4170 $Y=-1490
X1 1 2 3 ICV_6 $T=2920 0 0 0 $X=-1250 $Y=-1490
.ENDS
***************************************
.SUBCKT nmos_small
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_8
** N=4 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4
** N=4 EP=4 IP=8 FDC=1
M0 2 3 1 4 N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=9.8e-13 PD=2.98e-06 PS=2.98e-06 $X=-3310 $Y=-1325 $D=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4
** N=4 EP=4 IP=8 FDC=2
X0 1 2 3 4 ICV_9 $T=-1460 0 0 0 $X=-5460 $Y=-2800
X1 1 2 3 4 ICV_9 $T=0 0 0 0 $X=-4000 $Y=-2800
.ENDS
***************************************
.SUBCKT part1_2 A C B VSS OUT VDD
** N=8 EP=6 IP=71 FDC=39
X0 7 OUT C VDD ICV_3 $T=-3100 -4010 0 180 $X=-1090 $Y=-6295
X1 7 OUT C VDD ICV_3 $T=-180 -4010 0 180 $X=1830 $Y=-6295
X2 7 OUT C VDD ICV_3 $T=2740 -4010 0 180 $X=4750 $Y=-6295
X3 7 VDD B ICV_6 $T=8715 3900 0 0 $X=4545 $Y=2410
X4 7 VDD A ICV_7 $T=-15345 3900 0 0 $X=-19515 $Y=2410
X5 7 VDD A ICV_7 $T=-9505 3900 0 0 $X=-13675 $Y=2410
X6 7 VDD A ICV_7 $T=-3665 3900 0 0 $X=-7835 $Y=2410
X7 7 VDD B ICV_7 $T=2875 3900 0 0 $X=-1295 $Y=2410
X8 4 OUT A VSS ICV_9 $T=-22730 -4295 0 180 $X=-20290 $Y=-5720
X9 4 VSS B VSS ICV_9 $T=-13780 -4300 0 180 $X=-11340 $Y=-5725
X10 OUT VSS C VSS ICV_9 $T=-6380 -4295 0 180 $X=-3940 $Y=-5720
X11 4 OUT A VSS ICV_10 $T=-28570 -4295 0 180 $X=-26130 $Y=-5720
X12 4 OUT A VSS ICV_10 $T=-25650 -4295 0 180 $X=-23210 $Y=-5720
X13 4 VSS B VSS ICV_10 $T=-19620 -4300 0 180 $X=-17180 $Y=-5725
X14 4 VSS B VSS ICV_10 $T=-16700 -4300 0 180 $X=-14260 $Y=-5725
X15 OUT VSS C VSS ICV_10 $T=-12220 -4295 0 180 $X=-9780 $Y=-5720
X16 OUT VSS C VSS ICV_10 $T=-9300 -4295 0 180 $X=-6860 $Y=-5720
.ENDS
***************************************
