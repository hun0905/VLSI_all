* File: hw2_part2_2.pex.spi
* Created: Sun Nov 14 20:01:55 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw2_part2_2.pex.spi.pex"
.subckt hw2_part2_2  VDD VSS IN OUT1 OUT2 OUT3
* 
* OUT3	OUT3
* OUT2	OUT2
* OUT1	OUT1
* IN	IN
* VSS	VSS
* VDD	VDD
MM8 N_NET050_MM8_d N_NET062_MM8_g N_VSS_MM8_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.225e-12 AS=1.225e-12 PD=3.48e-06 PS=3.48e-06
MM9 N_NET054_MM9_d N_NET050_MM9_g N_VSS_MM9_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM9@5 N_NET054_MM9@5_d N_NET050_MM9@5_g N_VSS_MM9@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13 N_OUT1_MM13_d N_NET070_MM13_g N_VSS_MM13_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM9@4 N_NET054_MM9@4_d N_NET050_MM9@4_g N_VSS_MM9@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@25 N_OUT1_MM13@25_d N_NET070_MM13@25_g N_VSS_MM13@25_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM9@3 N_NET054_MM9@3_d N_NET050_MM9@3_g N_VSS_MM9@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@24 N_OUT1_MM13@24_d N_NET070_MM13@24_g N_VSS_MM13@24_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM9@2 N_NET054_MM9@2_d N_NET050_MM9@2_g N_VSS_MM9@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM13@23 N_OUT1_MM13@23_d N_NET070_MM13@23_g N_VSS_MM13@23_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@22 N_OUT1_MM13@22_d N_NET070_MM13@22_g N_VSS_MM13@22_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@21 N_OUT1_MM13@21_d N_NET070_MM13@21_g N_VSS_MM13@21_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11 N_NET0210_MM11_d N_NET054_MM11_g N_VSS_MM11_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM13@20 N_OUT1_MM13@20_d N_NET070_MM13@20_g N_VSS_MM13@20_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@25 N_NET0210_MM11@25_d N_NET054_MM11@25_g N_VSS_MM11@25_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@19 N_OUT1_MM13@19_d N_NET070_MM13@19_g N_VSS_MM13@19_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@24 N_NET0210_MM11@24_d N_NET054_MM11@24_g N_VSS_MM11@24_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@18 N_OUT1_MM13@18_d N_NET070_MM13@18_g N_VSS_MM13@18_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@23 N_NET0210_MM11@23_d N_NET054_MM11@23_g N_VSS_MM11@23_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@17 N_OUT1_MM13@17_d N_NET070_MM13@17_g N_VSS_MM13@17_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@22 N_NET0210_MM11@22_d N_NET054_MM11@22_g N_VSS_MM11@22_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@16 N_OUT1_MM13@16_d N_NET070_MM13@16_g N_VSS_MM13@16_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@21 N_NET0210_MM11@21_d N_NET054_MM11@21_g N_VSS_MM11@21_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@15 N_OUT1_MM13@15_d N_NET070_MM13@15_g N_VSS_MM13@15_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@20 N_NET0210_MM11@20_d N_NET054_MM11@20_g N_VSS_MM11@20_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@14 N_OUT1_MM13@14_d N_NET070_MM13@14_g N_VSS_MM13@14_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@19 N_NET0210_MM11@19_d N_NET054_MM11@19_g N_VSS_MM11@19_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@13 N_OUT1_MM13@13_d N_NET070_MM13@13_g N_VSS_MM13@13_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@18 N_NET0210_MM11@18_d N_NET054_MM11@18_g N_VSS_MM11@18_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@12 N_OUT1_MM13@12_d N_NET070_MM13@12_g N_VSS_MM13@12_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@17 N_NET0210_MM11@17_d N_NET054_MM11@17_g N_VSS_MM11@17_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@11 N_OUT1_MM13@11_d N_NET070_MM13@11_g N_VSS_MM13@11_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@16 N_NET0210_MM11@16_d N_NET054_MM11@16_g N_VSS_MM11@16_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@10 N_OUT1_MM13@10_d N_NET070_MM13@10_g N_VSS_MM13@10_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@15 N_NET0210_MM11@15_d N_NET054_MM11@15_g N_VSS_MM11@15_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@9 N_OUT1_MM13@9_d N_NET070_MM13@9_g N_VSS_MM13@9_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@14 N_NET0210_MM11@14_d N_NET054_MM11@14_g N_VSS_MM11@14_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@8 N_OUT1_MM13@8_d N_NET070_MM13@8_g N_VSS_MM13@8_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@13 N_NET0210_MM11@13_d N_NET054_MM11@13_g N_VSS_MM11@13_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@7 N_OUT1_MM13@7_d N_NET070_MM13@7_g N_VSS_MM13@7_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@12 N_NET0210_MM11@12_d N_NET054_MM11@12_g N_VSS_MM11@12_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@6 N_OUT1_MM13@6_d N_NET070_MM13@6_g N_VSS_MM13@6_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@11 N_NET0210_MM11@11_d N_NET054_MM11@11_g N_VSS_MM11@11_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@5 N_OUT1_MM13@5_d N_NET070_MM13@5_g N_VSS_MM13@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@10 N_NET0210_MM11@10_d N_NET054_MM11@10_g N_VSS_MM11@10_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@4 N_OUT1_MM13@4_d N_NET070_MM13@4_g N_VSS_MM13@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@9 N_NET0210_MM11@9_d N_NET054_MM11@9_g N_VSS_MM11@9_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@3 N_OUT1_MM13@3_d N_NET070_MM13@3_g N_VSS_MM13@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@8 N_NET0210_MM11@8_d N_NET054_MM11@8_g N_VSS_MM11@8_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM13@2 N_OUT1_MM13@2_d N_NET070_MM13@2_g N_VSS_MM13@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM11@7 N_NET0210_MM11@7_d N_NET054_MM11@7_g N_VSS_MM11@7_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@6 N_NET0210_MM11@6_d N_NET054_MM11@6_g N_VSS_MM11@6_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@5 N_NET0210_MM11@5_d N_NET054_MM11@5_g N_VSS_MM11@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@4 N_NET0210_MM11@4_d N_NET054_MM11@4_g N_VSS_MM11@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@3 N_NET0210_MM11@3_d N_NET054_MM11@3_g N_VSS_MM11@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@2 N_NET0210_MM11@2_d N_NET054_MM11@2_g N_VSS_MM11@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM22 N_NET0322_MM22_d N_NET074_MM22_g N_VSS_MM22_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM22@5 N_NET0322_MM22@5_d N_NET074_MM22@5_g N_VSS_MM22@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM22@4 N_NET0322_MM22@4_d N_NET074_MM22@4_g N_VSS_MM22@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM22@3 N_NET0322_MM22@3_d N_NET074_MM22@3_g N_VSS_MM22@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM22@2 N_NET0322_MM22@2_d N_NET074_MM22@2_g N_VSS_MM22@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM23 N_OUT2_MM23_d N_NET0322_MM23_g N_VSS_MM23_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM23@25 N_OUT2_MM23@25_d N_NET0322_MM23@25_g N_VSS_MM23@25_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@24 N_OUT2_MM23@24_d N_NET0322_MM23@24_g N_VSS_MM23@24_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@23 N_OUT2_MM23@23_d N_NET0322_MM23@23_g N_VSS_MM23@23_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@22 N_OUT2_MM23@22_d N_NET0322_MM23@22_g N_VSS_MM23@22_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM38 N_NET046_MM38_d N_NET0321_MM38_g N_VSS_MM38_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM23@21 N_OUT2_MM23@21_d N_NET0322_MM23@21_g N_VSS_MM23@21_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM38@5 N_NET046_MM38@5_d N_NET0321_MM38@5_g N_VSS_MM38@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@20 N_OUT2_MM23@20_d N_NET0322_MM23@20_g N_VSS_MM23@20_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM38@4 N_NET046_MM38@4_d N_NET0321_MM38@4_g N_VSS_MM38@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@19 N_OUT2_MM23@19_d N_NET0322_MM23@19_g N_VSS_MM23@19_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM38@3 N_NET046_MM38@3_d N_NET0321_MM38@3_g N_VSS_MM38@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@18 N_OUT2_MM23@18_d N_NET0322_MM23@18_g N_VSS_MM23@18_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM38@2 N_NET046_MM38@2_d N_NET0321_MM38@2_g N_VSS_MM38@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM23@17 N_OUT2_MM23@17_d N_NET0322_MM23@17_g N_VSS_MM23@17_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@16 N_OUT2_MM23@16_d N_NET0322_MM23@16_g N_VSS_MM23@16_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@15 N_OUT2_MM23@15_d N_NET0322_MM23@15_g N_VSS_MM23@15_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39 N_OUT3_MM39_d N_NET046_MM39_g N_VSS_MM39_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM23@14 N_OUT2_MM23@14_d N_NET0322_MM23@14_g N_VSS_MM23@14_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@25 N_OUT3_MM39@25_d N_NET046_MM39@25_g N_VSS_MM39@25_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@13 N_OUT2_MM23@13_d N_NET0322_MM23@13_g N_VSS_MM23@13_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@24 N_OUT3_MM39@24_d N_NET046_MM39@24_g N_VSS_MM39@24_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@12 N_OUT2_MM23@12_d N_NET0322_MM23@12_g N_VSS_MM23@12_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@23 N_OUT3_MM39@23_d N_NET046_MM39@23_g N_VSS_MM39@23_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@11 N_OUT2_MM23@11_d N_NET0322_MM23@11_g N_VSS_MM23@11_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@22 N_OUT3_MM39@22_d N_NET046_MM39@22_g N_VSS_MM39@22_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@10 N_OUT2_MM23@10_d N_NET0322_MM23@10_g N_VSS_MM23@10_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@21 N_OUT3_MM39@21_d N_NET046_MM39@21_g N_VSS_MM39@21_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@9 N_OUT2_MM23@9_d N_NET0322_MM23@9_g N_VSS_MM23@9_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@20 N_OUT3_MM39@20_d N_NET046_MM39@20_g N_VSS_MM39@20_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@8 N_OUT2_MM23@8_d N_NET0322_MM23@8_g N_VSS_MM23@8_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@19 N_OUT3_MM39@19_d N_NET046_MM39@19_g N_VSS_MM39@19_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@7 N_OUT2_MM23@7_d N_NET0322_MM23@7_g N_VSS_MM23@7_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@18 N_OUT3_MM39@18_d N_NET046_MM39@18_g N_VSS_MM39@18_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@6 N_OUT2_MM23@6_d N_NET0322_MM23@6_g N_VSS_MM23@6_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@17 N_OUT3_MM39@17_d N_NET046_MM39@17_g N_VSS_MM39@17_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@5 N_OUT2_MM23@5_d N_NET0322_MM23@5_g N_VSS_MM23@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@16 N_OUT3_MM39@16_d N_NET046_MM39@16_g N_VSS_MM39@16_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@4 N_OUT2_MM23@4_d N_NET0322_MM23@4_g N_VSS_MM23@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@15 N_OUT3_MM39@15_d N_NET046_MM39@15_g N_VSS_MM39@15_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@3 N_OUT2_MM23@3_d N_NET0322_MM23@3_g N_VSS_MM23@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@14 N_OUT3_MM39@14_d N_NET046_MM39@14_g N_VSS_MM39@14_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM23@2 N_OUT2_MM23@2_d N_NET0322_MM23@2_g N_VSS_MM23@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM39@13 N_OUT3_MM39@13_d N_NET046_MM39@13_g N_VSS_MM39@13_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@12 N_OUT3_MM39@12_d N_NET046_MM39@12_g N_VSS_MM39@12_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@11 N_OUT3_MM39@11_d N_NET046_MM39@11_g N_VSS_MM39@11_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@10 N_OUT3_MM39@10_d N_NET046_MM39@10_g N_VSS_MM39@10_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@9 N_OUT3_MM39@9_d N_NET046_MM39@9_g N_VSS_MM39@9_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@8 N_OUT3_MM39@8_d N_NET046_MM39@8_g N_VSS_MM39@8_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@7 N_OUT3_MM39@7_d N_NET046_MM39@7_g N_VSS_MM39@7_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@6 N_OUT3_MM39@6_d N_NET046_MM39@6_g N_VSS_MM39@6_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@5 N_OUT3_MM39@5_d N_NET046_MM39@5_g N_VSS_MM39@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@4 N_OUT3_MM39@4_d N_NET046_MM39@4_g N_VSS_MM39@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@3 N_OUT3_MM39@3_d N_NET046_MM39@3_g N_VSS_MM39@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM39@2 N_OUT3_MM39@2_d N_NET046_MM39@2_g N_VSS_MM39@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM10 N_NET058_MM10_d N_IN_MM10_g N_VSS_MM10_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM4 N_NET062_MM4_d N_NET058_MM4_g N_VSS_MM4_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM12 N_NET070_MM12_d N_NET0210_MM12_g N_VSS_MM12_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
MM12@5 N_NET070_MM12@5_d N_NET0210_MM12@5_g N_VSS_MM12@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
MM12@4 N_NET070_MM12@4_d N_NET0210_MM12@4_g N_VSS_MM12@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
MM12@3 N_NET070_MM12@3_d N_NET0210_MM12@3_g N_VSS_MM12@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
MM12@2 N_NET070_MM12@2_d N_NET0210_MM12@2_g N_VSS_MM12@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
MM26 N_NET090_MM26_d N_NET0210_MM26_g N_VSS_MM26_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM17 N_NET082_MM17_d N_NET0210_MM17_g N_VSS_MM17_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM27 N_NET0106_MM27_d N_NET090_MM27_g N_VSS_MM27_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM16 N_NET074_MM16_d N_NET082_MM16_g N_VSS_MM16_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM25 N_NET094_MM25_d N_NET0106_MM25_g N_VSS_MM25_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM24 N_NET098_MM24_d N_NET094_MM24_g N_VSS_MM24_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM37 N_NET0323_MM37_d N_NET098_MM37_g N_VSS_MM37_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM36 N_NET0321_MM36_d N_NET0323_MM36_g N_VSS_MM36_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM15 N_OUT1_MM15_d N_NET070_MM15_g N_VDD_MM15_s N_VDD_MM14@3_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM15@25 N_OUT1_MM15@25_d N_NET070_MM15@25_g N_VDD_MM15@25_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@24 N_OUT1_MM15@24_d N_NET070_MM15@24_g N_VDD_MM15@24_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@23 N_OUT1_MM15@23_d N_NET070_MM15@23_g N_VDD_MM15@23_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@22 N_OUT1_MM15@22_d N_NET070_MM15@22_g N_VDD_MM15@22_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@21 N_OUT1_MM15@21_d N_NET070_MM15@21_g N_VDD_MM15@21_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7 N_NET0210_MM7_d N_NET054_MM7_g N_VDD_MM7_s N_VDD_MM5@3_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM15@20 N_OUT1_MM15@20_d N_NET070_MM15@20_g N_VDD_MM15@20_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@25 N_NET0210_MM7@25_d N_NET054_MM7@25_g N_VDD_MM7@25_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@19 N_OUT1_MM15@19_d N_NET070_MM15@19_g N_VDD_MM15@19_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@24 N_NET0210_MM7@24_d N_NET054_MM7@24_g N_VDD_MM7@24_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@18 N_OUT1_MM15@18_d N_NET070_MM15@18_g N_VDD_MM15@18_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@23 N_NET0210_MM7@23_d N_NET054_MM7@23_g N_VDD_MM7@23_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@17 N_OUT1_MM15@17_d N_NET070_MM15@17_g N_VDD_MM15@17_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@22 N_NET0210_MM7@22_d N_NET054_MM7@22_g N_VDD_MM7@22_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@16 N_OUT1_MM15@16_d N_NET070_MM15@16_g N_VDD_MM15@16_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@21 N_NET0210_MM7@21_d N_NET054_MM7@21_g N_VDD_MM7@21_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@15 N_OUT1_MM15@15_d N_NET070_MM15@15_g N_VDD_MM15@15_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@20 N_NET0210_MM7@20_d N_NET054_MM7@20_g N_VDD_MM7@20_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@14 N_OUT1_MM15@14_d N_NET070_MM15@14_g N_VDD_MM15@14_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@19 N_NET0210_MM7@19_d N_NET054_MM7@19_g N_VDD_MM7@19_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@13 N_OUT1_MM15@13_d N_NET070_MM15@13_g N_VDD_MM15@13_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@18 N_NET0210_MM7@18_d N_NET054_MM7@18_g N_VDD_MM7@18_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@12 N_OUT1_MM15@12_d N_NET070_MM15@12_g N_VDD_MM15@12_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@17 N_NET0210_MM7@17_d N_NET054_MM7@17_g N_VDD_MM7@17_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@11 N_OUT1_MM15@11_d N_NET070_MM15@11_g N_VDD_MM15@11_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@16 N_NET0210_MM7@16_d N_NET054_MM7@16_g N_VDD_MM7@16_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@10 N_OUT1_MM15@10_d N_NET070_MM15@10_g N_VDD_MM15@10_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@15 N_NET0210_MM7@15_d N_NET054_MM7@15_g N_VDD_MM7@15_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@9 N_OUT1_MM15@9_d N_NET070_MM15@9_g N_VDD_MM15@9_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@14 N_NET0210_MM7@14_d N_NET054_MM7@14_g N_VDD_MM7@14_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@8 N_OUT1_MM15@8_d N_NET070_MM15@8_g N_VDD_MM15@8_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@13 N_NET0210_MM7@13_d N_NET054_MM7@13_g N_VDD_MM7@13_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@7 N_OUT1_MM15@7_d N_NET070_MM15@7_g N_VDD_MM15@7_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@12 N_NET0210_MM7@12_d N_NET054_MM7@12_g N_VDD_MM7@12_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@6 N_OUT1_MM15@6_d N_NET070_MM15@6_g N_VDD_MM15@6_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@11 N_NET0210_MM7@11_d N_NET054_MM7@11_g N_VDD_MM7@11_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@5 N_OUT1_MM15@5_d N_NET070_MM15@5_g N_VDD_MM15@5_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@10 N_NET0210_MM7@10_d N_NET054_MM7@10_g N_VDD_MM7@10_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@4 N_OUT1_MM15@4_d N_NET070_MM15@4_g N_VDD_MM15@4_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@9 N_NET0210_MM7@9_d N_NET054_MM7@9_g N_VDD_MM7@9_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@3 N_OUT1_MM15@3_d N_NET070_MM15@3_g N_VDD_MM15@3_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@8 N_NET0210_MM7@8_d N_NET054_MM7@8_g N_VDD_MM7@8_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM15@2 N_OUT1_MM15@2_d N_NET070_MM15@2_g N_VDD_MM15@2_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM7@7 N_NET0210_MM7@7_d N_NET054_MM7@7_g N_VDD_MM7@7_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@6 N_NET0210_MM7@6_d N_NET054_MM7@6_g N_VDD_MM7@6_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@5 N_NET0210_MM7@5_d N_NET054_MM7@5_g N_VDD_MM7@5_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@4 N_NET0210_MM7@4_d N_NET054_MM7@4_g N_VDD_MM7@4_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@3 N_NET0210_MM7@3_d N_NET054_MM7@3_g N_VDD_MM7@3_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@2 N_NET0210_MM7@2_d N_NET054_MM7@2_g N_VDD_MM7@2_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM21 N_OUT2_MM21_d N_NET0322_MM21_g N_VDD_MM21_s N_VDD_MM20@3_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM21@25 N_OUT2_MM21@25_d N_NET0322_MM21@25_g N_VDD_MM21@25_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@24 N_OUT2_MM21@24_d N_NET0322_MM21@24_g N_VDD_MM21@24_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@23 N_OUT2_MM21@23_d N_NET0322_MM21@23_g N_VDD_MM21@23_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@22 N_OUT2_MM21@22_d N_NET0322_MM21@22_g N_VDD_MM21@22_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@21 N_OUT2_MM21@21_d N_NET0322_MM21@21_g N_VDD_MM21@21_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@20 N_OUT2_MM21@20_d N_NET0322_MM21@20_g N_VDD_MM21@20_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@19 N_OUT2_MM21@19_d N_NET0322_MM21@19_g N_VDD_MM21@19_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@18 N_OUT2_MM21@18_d N_NET0322_MM21@18_g N_VDD_MM21@18_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@17 N_OUT2_MM21@17_d N_NET0322_MM21@17_g N_VDD_MM21@17_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@16 N_OUT2_MM21@16_d N_NET0322_MM21@16_g N_VDD_MM21@16_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@15 N_OUT2_MM21@15_d N_NET0322_MM21@15_g N_VDD_MM21@15_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35 N_OUT3_MM35_d N_NET046_MM35_g N_VDD_MM35_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM21@14 N_OUT2_MM21@14_d N_NET0322_MM21@14_g N_VDD_MM21@14_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@25 N_OUT3_MM35@25_d N_NET046_MM35@25_g N_VDD_MM35@25_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@13 N_OUT2_MM21@13_d N_NET0322_MM21@13_g N_VDD_MM21@13_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@24 N_OUT3_MM35@24_d N_NET046_MM35@24_g N_VDD_MM35@24_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@12 N_OUT2_MM21@12_d N_NET0322_MM21@12_g N_VDD_MM21@12_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@23 N_OUT3_MM35@23_d N_NET046_MM35@23_g N_VDD_MM35@23_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@11 N_OUT2_MM21@11_d N_NET0322_MM21@11_g N_VDD_MM21@11_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@22 N_OUT3_MM35@22_d N_NET046_MM35@22_g N_VDD_MM35@22_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@10 N_OUT2_MM21@10_d N_NET0322_MM21@10_g N_VDD_MM21@10_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@21 N_OUT3_MM35@21_d N_NET046_MM35@21_g N_VDD_MM35@21_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@9 N_OUT2_MM21@9_d N_NET0322_MM21@9_g N_VDD_MM21@9_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@20 N_OUT3_MM35@20_d N_NET046_MM35@20_g N_VDD_MM35@20_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@8 N_OUT2_MM21@8_d N_NET0322_MM21@8_g N_VDD_MM21@8_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@19 N_OUT3_MM35@19_d N_NET046_MM35@19_g N_VDD_MM35@19_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@7 N_OUT2_MM21@7_d N_NET0322_MM21@7_g N_VDD_MM21@7_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@18 N_OUT3_MM35@18_d N_NET046_MM35@18_g N_VDD_MM35@18_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@6 N_OUT2_MM21@6_d N_NET0322_MM21@6_g N_VDD_MM21@6_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@17 N_OUT3_MM35@17_d N_NET046_MM35@17_g N_VDD_MM35@17_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@5 N_OUT2_MM21@5_d N_NET0322_MM21@5_g N_VDD_MM21@5_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@16 N_OUT3_MM35@16_d N_NET046_MM35@16_g N_VDD_MM35@16_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@4 N_OUT2_MM21@4_d N_NET0322_MM21@4_g N_VDD_MM21@4_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@15 N_OUT3_MM35@15_d N_NET046_MM35@15_g N_VDD_MM35@15_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@3 N_OUT2_MM21@3_d N_NET0322_MM21@3_g N_VDD_MM21@3_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@14 N_OUT3_MM35@14_d N_NET046_MM35@14_g N_VDD_MM35@14_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM21@2 N_OUT2_MM21@2_d N_NET0322_MM21@2_g N_VDD_MM21@2_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM35@13 N_OUT3_MM35@13_d N_NET046_MM35@13_g N_VDD_MM35@13_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@12 N_OUT3_MM35@12_d N_NET046_MM35@12_g N_VDD_MM35@12_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@11 N_OUT3_MM35@11_d N_NET046_MM35@11_g N_VDD_MM35@11_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@10 N_OUT3_MM35@10_d N_NET046_MM35@10_g N_VDD_MM35@10_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@9 N_OUT3_MM35@9_d N_NET046_MM35@9_g N_VDD_MM35@9_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@8 N_OUT3_MM35@8_d N_NET046_MM35@8_g N_VDD_MM35@8_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@7 N_OUT3_MM35@7_d N_NET046_MM35@7_g N_VDD_MM35@7_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@6 N_OUT3_MM35@6_d N_NET046_MM35@6_g N_VDD_MM35@6_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@5 N_OUT3_MM35@5_d N_NET046_MM35@5_g N_VDD_MM35@5_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@4 N_OUT3_MM35@4_d N_NET046_MM35@4_g N_VDD_MM35@4_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@3 N_OUT3_MM35@3_d N_NET046_MM35@3_g N_VDD_MM35@3_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM35@2 N_OUT3_MM35@2_d N_NET046_MM35@2_g N_VDD_MM35@2_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM3 N_NET050_MM3_d N_NET062_MM3_g N_VDD_MM3_s N_VDD_MM5@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM14 N_NET070_MM14_d N_NET0210_MM14_g N_VDD_MM14_s N_VDD_MM14@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=4.7175e-13 PD=2.83e-06 PS=5.1e-07
MM5 N_NET054_MM5_d N_NET050_MM5_g N_VDD_MM5_s N_VDD_MM5@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=4.7175e-13 PD=2.83e-06 PS=5.1e-07
MM20 N_NET0322_MM20_d N_NET074_MM20_g N_VDD_MM20_s N_VDD_MM20@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=4.7175e-13 PD=2.83e-06 PS=5.1e-07
MM34 N_NET046_MM34_d N_NET0321_MM34_g N_VDD_MM34_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=4.7175e-13 PD=2.83e-06 PS=5.1e-07
MM14@5 N_NET070_MM14@5_d N_NET0210_MM14@5_g N_VDD_MM14@5_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
MM14@4 N_NET070_MM14@4_d N_NET0210_MM14@4_g N_VDD_MM14@4_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM5@5 N_NET054_MM5@5_d N_NET050_MM5@5_g N_VDD_MM5@5_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
MM5@4 N_NET054_MM5@4_d N_NET050_MM5@4_g N_VDD_MM5@4_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM20@5 N_NET0322_MM20@5_d N_NET074_MM20@5_g N_VDD_MM20@5_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
MM20@4 N_NET0322_MM20@4_d N_NET074_MM20@4_g N_VDD_MM20@4_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM34@5 N_NET046_MM34@5_d N_NET0321_MM34@5_g N_VDD_MM34@5_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
MM34@4 N_NET046_MM34@4_d N_NET0321_MM34@4_g N_VDD_MM34@4_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM14@3 N_NET070_MM14@3_d N_NET0210_MM14@3_g N_VDD_MM14@3_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM14@2 N_NET070_MM14@2_d N_NET0210_MM14@2_g N_VDD_MM14@2_s N_VDD_MM14@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM5@3 N_NET054_MM5@3_d N_NET050_MM5@3_g N_VDD_MM5@3_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM5@2 N_NET054_MM5@2_d N_NET050_MM5@2_g N_VDD_MM5@2_s N_VDD_MM5@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM20@3 N_NET0322_MM20@3_d N_NET074_MM20@3_g N_VDD_MM20@3_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM20@2 N_NET0322_MM20@2_d N_NET074_MM20@2_g N_VDD_MM20@2_s N_VDD_MM20@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM34@3 N_NET046_MM34@3_d N_NET0321_MM34@3_g N_VDD_MM34@3_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM34@2 N_NET046_MM34@2_d N_NET0321_MM34@2_g N_VDD_MM34@2_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM6 N_NET058_MM6_d N_IN_MM6_g N_VDD_MM6_s N_VDD_MM5@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM0 N_NET062_MM0_d N_NET058_MM0_g N_VDD_MM0_s N_VDD_MM5@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM30 N_NET090_MM30_d N_NET0210_MM30_g N_VDD_MM30_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM31 N_NET0106_MM31_d N_NET090_MM31_g N_VDD_MM31_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM19 N_NET082_MM19_d N_NET0210_MM19_g N_VDD_MM19_s N_VDD_MM20@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM18 N_NET074_MM18_d N_NET082_MM18_g N_VDD_MM18_s N_VDD_MM20@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM29 N_NET094_MM29_d N_NET0106_MM29_g N_VDD_MM29_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM28 N_NET098_MM28_d N_NET094_MM28_g N_VDD_MM28_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM33 N_NET0323_MM33_d N_NET098_MM33_g N_VDD_MM33_s N_VDD_MM34@3_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM32 N_NET0321_MM32_d N_NET0323_MM32_g N_VDD_MM32_s N_VDD_MM34@3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
*
.include "hw2_part2_2.pex.spi.HW2_PART2_2.pxi"
*
.ends
*
*
