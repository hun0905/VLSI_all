* File: hw2_part1_2.pex.spi
* Created: Thu Nov 11 10:56:45 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw2_part1_2.pex.spi.pex"
.subckt hw2_part1_2  VSS A B VDD C OUT
* 
* OUT	OUT
* C	C
* VDD	VDD
* B	B
* A	A
* VSS	VSS
MM3 N_OUT_MM3_d N_A_MM3_g N_noxref_4_MM3_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06
MM3@5 N_OUT_MM3@5_d N_A_MM3@5_g N_noxref_4_MM3@5_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM3@4 N_OUT_MM3@4_d N_A_MM3@4_g N_noxref_4_MM3@4_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM3@3 N_OUT_MM3@3_d N_A_MM3@3_g N_noxref_4_MM3@3_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM3@2 N_OUT_MM3@2_d N_A_MM3@2_g N_noxref_4_MM3@2_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07
MM4 N_noxref_4_MM4_d N_B_MM4_g N_VSS_MM4_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07
MM4@5 N_noxref_4_MM4@5_d N_B_MM4@5_g N_VSS_MM4@5_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM4@4 N_noxref_4_MM4@4_d N_B_MM4@4_g N_VSS_MM4@4_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM4@3 N_noxref_4_MM4@3_d N_B_MM4@3_g N_VSS_MM4@3_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM4@2 N_noxref_4_MM4@2_d N_B_MM4@2_g N_VSS_MM4@2_s N_VSS_MM3_b N_18 L=1.8e-07
+ W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06
MM5 N_OUT_MM5_d N_C_MM5_g N_VSS_MM5_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07
MM5@5 N_OUT_MM5@5_d N_C_MM5@5_g N_VSS_MM5@5_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM5@4 N_OUT_MM5@4_d N_C_MM5@4_g N_VSS_MM5@4_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM5@3 N_OUT_MM5@3_d N_C_MM5@3_g N_VSS_MM5@3_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07
MM5@2 N_OUT_MM5@2_d N_C_MM5@2_g N_VSS_MM5@2_s N_VSS_MM3_b N_18 L=1.8e-07 W=2e-06
+ AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06
MM0 N_noxref_8_MM0_d N_A_MM0_g N_VDD_MM0_s N_VDD_MM0_b P_18 L=1.8e-07 W=2.5e-06
+ AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM0@12 N_noxref_8_MM0@12_d N_A_MM0@12_g N_VDD_MM0@12_s N_VDD_MM0_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@11 N_noxref_8_MM0@11_d N_A_MM0@11_g N_VDD_MM0@11_s N_VDD_MM0_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@10 N_noxref_8_MM0@10_d N_A_MM0@10_g N_VDD_MM0@10_s N_VDD_MM0_b P_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@9 N_noxref_8_MM0@9_d N_A_MM0@9_g N_VDD_MM0@9_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@8 N_noxref_8_MM0@8_d N_A_MM0@8_g N_VDD_MM0@8_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@7 N_noxref_8_MM0@7_d N_A_MM0@7_g N_VDD_MM0@7_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@6 N_noxref_8_MM0@6_d N_A_MM0@6_g N_VDD_MM0@6_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@5 N_noxref_8_MM0@5_d N_A_MM0@5_g N_VDD_MM0@5_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@4 N_noxref_8_MM0@4_d N_A_MM0@4_g N_VDD_MM0@4_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@3 N_noxref_8_MM0@3_d N_A_MM0@3_g N_VDD_MM0@3_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM0@2 N_noxref_8_MM0@2_d N_A_MM0@2_g N_VDD_MM0@2_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM1 N_noxref_8_MM1_d N_B_MM1_g N_VDD_MM1_s N_VDD_MM0_b P_18 L=1.8e-07 W=2.5e-06
+ AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM1@6 N_noxref_8_MM1@6_d N_B_MM1@6_g N_VDD_MM1@6_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM1@5 N_noxref_8_MM1@5_d N_B_MM1@5_g N_VDD_MM1@5_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM1@4 N_noxref_8_MM1@4_d N_B_MM1@4_g N_VDD_MM1@4_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM1@3 N_noxref_8_MM1@3_d N_B_MM1@3_g N_VDD_MM1@3_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM1@2 N_noxref_8_MM1@2_d N_B_MM1@2_g N_VDD_MM1@2_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM2 N_OUT_MM2_d N_C_MM2_g N_noxref_8_MM2_s N_VDD_MM0_b P_18 L=1.8e-07 W=2.5e-06
+ AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM2@6 N_OUT_MM2@6_d N_C_MM2@6_g N_noxref_8_MM2@6_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM2@5 N_OUT_MM2@5_d N_C_MM2@5_g N_noxref_8_MM2@5_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM2@4 N_OUT_MM2@4_d N_C_MM2@4_g N_noxref_8_MM2@4_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM2@3 N_OUT_MM2@3_d N_C_MM2@3_g N_noxref_8_MM2@3_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM2@2 N_OUT_MM2@2_d N_C_MM2@2_g N_noxref_8_MM2@2_s N_VDD_MM0_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
*
.include "hw2_part1_2.pex.spi.HW2_PART1_2.pxi"
*
.ends
*
*
