************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: and
* View Name:     schematic
* Netlisted on:  Jan 16 10:06:55 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    and
* View Name:    schematic
************************************************************************

.SUBCKT and A B OUT VDD VSS
*.PININFO A:I B:I OUT:O VDD:B VSS:B
MM10 OUT net067 VSS VSS N_18 W=500.0n L=180.00n m=1
MM5 net44 B VSS VSS N_18 W=500.0n L=180.00n m=1
MM4 net067 A net44 VSS N_18 W=500.0n L=180.00n m=1
MM9 OUT net067 VDD VDD P_18 W=500.0n L=180.00n m=3
MM1 net067 A VDD VDD P_18 W=500.0n L=180.00n m=3
MM0 net067 B VDD VDD P_18 W=500.0n L=180.00n m=3
.ENDS

