* File: Final_all_v1.pex.spi
* Created: Mon Jan 17 03:41:12 2022
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "Final_all_v1.pex.spi.pex"
.subckt Final  YOUT<0> YOUT<1> YOUT<2> YOUT<3> YOUT<4> YOUT<5> YOUT<6> YOUT<7>
+ DOUT<0> SO<0> DOUT<1> SO<1> VDD CLK WLEN VSS SAEN BL<0> BL<1> BL<2> BL<3>
+ BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15>
+ X_SEL<5> X_SEL<2> X_SEL<4> X_SEL<1> X_SEL<3> X_SEL<0> WL<63> WL<62> WL<61>
+ WL<60> WL<59> WL<58> WL<57> WL<56> WL<55> WL<54> WL<53> WL<52> WL<51> WL<50>
+ WL<49> WL<48> WL<47> WL<46> WL<45> WL<44> WL<43> WL<42> WL<41> WL<40> WL<39>
+ WL<38> WL<37> WL<36> WL<35> WL<34> WL<33> WL<32> WL<31> WL<30> WL<29> WL<28>
+ WL<27> WL<26> WL<25> WL<24> WL<23> WL<22> WL<21> WL<20> WL<19> WL<18> WL<17>
+ WL<16> WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> WL<9> WL<8> WL<7> WL<6> WL<5>
+ WL<4> WL<3> WL<2> WL<1> WL<0> DL<0> DL<1> Y_SEL<0> Y_SEL<2> Y_SEL<1> VREF A<2>
+ A<1> A<0> A<6> A<7> A<8> A<3> A<4> A<5>
* 
* A<5>	A<5>
* A<4>	A<4>
* A<3>	A<3>
* A<8>	A<8>
* A<7>	A<7>
* A<6>	A<6>
* A<0>	A<0>
* A<1>	A<1>
* A<2>	A<2>
* VREF	VREF
* Y_SEL<1>	Y_SEL<1>
* Y_SEL<2>	Y_SEL<2>
* Y_SEL<0>	Y_SEL<0>
* DL<1>	DL<1>
* DL<0>	DL<0>
* WL<0>	WL<0>
* WL<1>	WL<1>
* WL<2>	WL<2>
* WL<3>	WL<3>
* WL<4>	WL<4>
* WL<5>	WL<5>
* WL<6>	WL<6>
* WL<7>	WL<7>
* WL<8>	WL<8>
* WL<9>	WL<9>
* WL<10>	WL<10>
* WL<11>	WL<11>
* WL<12>	WL<12>
* WL<13>	WL<13>
* WL<14>	WL<14>
* WL<15>	WL<15>
* WL<16>	WL<16>
* WL<17>	WL<17>
* WL<18>	WL<18>
* WL<19>	WL<19>
* WL<20>	WL<20>
* WL<21>	WL<21>
* WL<22>	WL<22>
* WL<23>	WL<23>
* WL<24>	WL<24>
* WL<25>	WL<25>
* WL<26>	WL<26>
* WL<27>	WL<27>
* WL<28>	WL<28>
* WL<29>	WL<29>
* WL<30>	WL<30>
* WL<31>	WL<31>
* WL<32>	WL<32>
* WL<33>	WL<33>
* WL<34>	WL<34>
* WL<35>	WL<35>
* WL<36>	WL<36>
* WL<37>	WL<37>
* WL<38>	WL<38>
* WL<39>	WL<39>
* WL<40>	WL<40>
* WL<41>	WL<41>
* WL<42>	WL<42>
* WL<43>	WL<43>
* WL<44>	WL<44>
* WL<45>	WL<45>
* WL<46>	WL<46>
* WL<47>	WL<47>
* WL<48>	WL<48>
* WL<49>	WL<49>
* WL<50>	WL<50>
* WL<51>	WL<51>
* WL<52>	WL<52>
* WL<53>	WL<53>
* WL<54>	WL<54>
* WL<55>	WL<55>
* WL<56>	WL<56>
* WL<57>	WL<57>
* WL<58>	WL<58>
* WL<59>	WL<59>
* WL<60>	WL<60>
* WL<61>	WL<61>
* WL<62>	WL<62>
* WL<63>	WL<63>
* X_SEL<0>	X_SEL<0>
* X_SEL<3>	X_SEL<3>
* X_SEL<1>	X_SEL<1>
* X_SEL<4>	X_SEL<4>
* X_SEL<2>	X_SEL<2>
* X_SEL<5>	X_SEL<5>
* BL<15>	BL<15>
* BL<14>	BL<14>
* BL<13>	BL<13>
* BL<12>	BL<12>
* BL<11>	BL<11>
* BL<10>	BL<10>
* BL<9>	BL<9>
* BL<8>	BL<8>
* BL<7>	BL<7>
* BL<6>	BL<6>
* BL<5>	BL<5>
* BL<4>	BL<4>
* BL<3>	BL<3>
* BL<2>	BL<2>
* BL<1>	BL<1>
* BL<0>	BL<0>
* SAEN	SAEN
* VSS	VSS
* WL_EN	WL_EN
* CLK	CLK
* VDD	VDD
* SO<1>	SO<1>
* DOUT<1>	DOUT<1>
* SO<0>	SO<0>
* DOUT<0>	DOUT<0>
* YOUT<7>	YOUT<7>
* YOUT<6>	YOUT<6>
* YOUT<5>	YOUT<5>
* YOUT<4>	YOUT<4>
* YOUT<3>	YOUT<3>
* YOUT<2>	YOUT<2>
* YOUT<1>	YOUT<1>
* YOUT<0>	YOUT<0>
mXI9/XI0/XI10/MM10 N_XI9/XI0/NET0116_XI9/XI0/XI10/MM10_d
+ N_X_SEL<3>_XI9/XI0/XI10/MM10_g N_VSS_XI9/XI0/XI10/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI9/XI0/XI11/MM10 N_XI9/XI0/NET0105_XI9/XI0/XI11/MM10_d
+ N_X_SEL<4>_XI9/XI0/XI11/MM10_g N_VSS_XI9/XI0/XI11/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI9/XI0/XI8/MM10 N_XI9/XI0/NET0158_XI9/XI0/XI8/MM10_d
+ N_X_SEL<5>_XI9/XI0/XI8/MM10_g N_VSS_XI9/XI0/XI8/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI9/XI1/XI10/MM10 N_XI9/XI1/NET0116_XI9/XI1/XI10/MM10_d
+ N_X_SEL<0>_XI9/XI1/XI10/MM10_g N_VSS_XI9/XI1/XI10/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI9/XI1/XI11/MM10 N_XI9/XI1/NET0105_XI9/XI1/XI11/MM10_d
+ N_X_SEL<1>_XI9/XI1/XI11/MM10_g N_VSS_XI9/XI1/XI11/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI9/XI1/XI8/MM10 N_XI9/XI1/NET0158_XI9/XI1/XI8/MM10_d
+ N_X_SEL<2>_XI9/XI1/XI8/MM10_g N_VSS_XI9/XI1/XI8/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI9/XI0/XI7/MM11 N_XI9/XI0/XI7/NET030_XI9/XI0/XI7/MM11_d
+ N_WLEN_XI9/XI0/XI7/MM11_g N_VSS_XI9/XI0/XI7/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI7/MM6 N_XI9/XI0/XI7/NET40_XI9/XI0/XI7/MM6_d
+ N_X_SEL<3>_XI9/XI0/XI7/MM6_g N_XI9/XI0/XI7/NET030_XI9/XI0/XI7/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI7/MM5 N_XI9/XI0/XI7/NET44_XI9/XI0/XI7/MM5_d
+ N_X_SEL<4>_XI9/XI0/XI7/MM5_g N_XI9/XI0/XI7/NET40_XI9/XI0/XI7/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI7/MM4 N_XI9/NET17_XI9/XI0/XI7/MM4_d N_X_SEL<5>_XI9/XI0/XI7/MM4_g
+ N_XI9/XI0/XI7/NET44_XI9/XI0/XI7/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI6/MM11 N_XI9/XI0/XI6/NET030_XI9/XI0/XI6/MM11_d
+ N_WLEN_XI9/XI0/XI6/MM11_g N_VSS_XI9/XI0/XI6/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI6/MM6 N_XI9/XI0/XI6/NET40_XI9/XI0/XI6/MM6_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI6/MM6_g N_XI9/XI0/XI6/NET030_XI9/XI0/XI6/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI6/MM5 N_XI9/XI0/XI6/NET44_XI9/XI0/XI6/MM5_d
+ N_X_SEL<4>_XI9/XI0/XI6/MM5_g N_XI9/XI0/XI6/NET40_XI9/XI0/XI6/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI6/MM4 N_XI9/NET18_XI9/XI0/XI6/MM4_d N_X_SEL<5>_XI9/XI0/XI6/MM4_g
+ N_XI9/XI0/XI6/NET44_XI9/XI0/XI6/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI5/MM11 N_XI9/XI0/XI5/NET030_XI9/XI0/XI5/MM11_d
+ N_WLEN_XI9/XI0/XI5/MM11_g N_VSS_XI9/XI0/XI5/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI5/MM6 N_XI9/XI0/XI5/NET40_XI9/XI0/XI5/MM6_d
+ N_X_SEL<3>_XI9/XI0/XI5/MM6_g N_XI9/XI0/XI5/NET030_XI9/XI0/XI5/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI5/MM5 N_XI9/XI0/XI5/NET44_XI9/XI0/XI5/MM5_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI5/MM5_g N_XI9/XI0/XI5/NET40_XI9/XI0/XI5/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI5/MM4 N_XI9/NET19_XI9/XI0/XI5/MM4_d N_X_SEL<5>_XI9/XI0/XI5/MM4_g
+ N_XI9/XI0/XI5/NET44_XI9/XI0/XI5/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI4/MM11 N_XI9/XI0/XI4/NET030_XI9/XI0/XI4/MM11_d
+ N_WLEN_XI9/XI0/XI4/MM11_g N_VSS_XI9/XI0/XI4/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI4/MM6 N_XI9/XI0/XI4/NET40_XI9/XI0/XI4/MM6_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI4/MM6_g N_XI9/XI0/XI4/NET030_XI9/XI0/XI4/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI4/MM5 N_XI9/XI0/XI4/NET44_XI9/XI0/XI4/MM5_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI4/MM5_g N_XI9/XI0/XI4/NET40_XI9/XI0/XI4/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI4/MM4 N_XI9/NET20_XI9/XI0/XI4/MM4_d N_X_SEL<5>_XI9/XI0/XI4/MM4_g
+ N_XI9/XI0/XI4/NET44_XI9/XI0/XI4/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI3/MM11 N_XI9/XI0/XI3/NET030_XI9/XI0/XI3/MM11_d
+ N_WLEN_XI9/XI0/XI3/MM11_g N_VSS_XI9/XI0/XI3/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI3/MM6 N_XI9/XI0/XI3/NET40_XI9/XI0/XI3/MM6_d
+ N_X_SEL<3>_XI9/XI0/XI3/MM6_g N_XI9/XI0/XI3/NET030_XI9/XI0/XI3/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI3/MM5 N_XI9/XI0/XI3/NET44_XI9/XI0/XI3/MM5_d
+ N_X_SEL<4>_XI9/XI0/XI3/MM5_g N_XI9/XI0/XI3/NET40_XI9/XI0/XI3/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI3/MM4 N_XI9/NET21_XI9/XI0/XI3/MM4_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI3/MM4_g N_XI9/XI0/XI3/NET44_XI9/XI0/XI3/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI2/MM11 N_XI9/XI0/XI2/NET030_XI9/XI0/XI2/MM11_d
+ N_WLEN_XI9/XI0/XI2/MM11_g N_VSS_XI9/XI0/XI2/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI2/MM6 N_XI9/XI0/XI2/NET40_XI9/XI0/XI2/MM6_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI2/MM6_g N_XI9/XI0/XI2/NET030_XI9/XI0/XI2/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI2/MM5 N_XI9/XI0/XI2/NET44_XI9/XI0/XI2/MM5_d
+ N_X_SEL<4>_XI9/XI0/XI2/MM5_g N_XI9/XI0/XI2/NET40_XI9/XI0/XI2/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI2/MM4 N_XI9/NET22_XI9/XI0/XI2/MM4_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI2/MM4_g N_XI9/XI0/XI2/NET44_XI9/XI0/XI2/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI1/MM11 N_XI9/XI0/XI1/NET030_XI9/XI0/XI1/MM11_d
+ N_WLEN_XI9/XI0/XI1/MM11_g N_VSS_XI9/XI0/XI1/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI1/MM6 N_XI9/XI0/XI1/NET40_XI9/XI0/XI1/MM6_d
+ N_X_SEL<3>_XI9/XI0/XI1/MM6_g N_XI9/XI0/XI1/NET030_XI9/XI0/XI1/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI1/MM5 N_XI9/XI0/XI1/NET44_XI9/XI0/XI1/MM5_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI1/MM5_g N_XI9/XI0/XI1/NET40_XI9/XI0/XI1/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI1/MM4 N_XI9/NET23_XI9/XI0/XI1/MM4_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI1/MM4_g N_XI9/XI0/XI1/NET44_XI9/XI0/XI1/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI0/MM11 N_XI9/XI0/XI0/NET030_XI9/XI0/XI0/MM11_d
+ N_WLEN_XI9/XI0/XI0/MM11_g N_VSS_XI9/XI0/XI0/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI0/XI0/MM6 N_XI9/XI0/XI0/NET40_XI9/XI0/XI0/MM6_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI0/MM6_g N_XI9/XI0/XI0/NET030_XI9/XI0/XI0/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI0/MM5 N_XI9/XI0/XI0/NET44_XI9/XI0/XI0/MM5_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI0/MM5_g N_XI9/XI0/XI0/NET40_XI9/XI0/XI0/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI0/XI0/MM4 N_XI9/NET24_XI9/XI0/XI0/MM4_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI0/MM4_g N_XI9/XI0/XI0/NET44_XI9/XI0/XI0/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI7/MM11 N_XI9/XI1/XI7/NET030_XI9/XI1/XI7/MM11_d
+ N_WLEN_XI9/XI1/XI7/MM11_g N_VSS_XI9/XI1/XI7/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI7/MM6 N_XI9/XI1/XI7/NET40_XI9/XI1/XI7/MM6_d
+ N_X_SEL<0>_XI9/XI1/XI7/MM6_g N_XI9/XI1/XI7/NET030_XI9/XI1/XI7/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI7/MM5 N_XI9/XI1/XI7/NET44_XI9/XI1/XI7/MM5_d
+ N_X_SEL<1>_XI9/XI1/XI7/MM5_g N_XI9/XI1/XI7/NET40_XI9/XI1/XI7/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI7/MM4 N_XI9/NET4_XI9/XI1/XI7/MM4_d N_X_SEL<2>_XI9/XI1/XI7/MM4_g
+ N_XI9/XI1/XI7/NET44_XI9/XI1/XI7/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI6/MM11 N_XI9/XI1/XI6/NET030_XI9/XI1/XI6/MM11_d
+ N_WLEN_XI9/XI1/XI6/MM11_g N_VSS_XI9/XI1/XI6/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI6/MM6 N_XI9/XI1/XI6/NET40_XI9/XI1/XI6/MM6_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI6/MM6_g N_XI9/XI1/XI6/NET030_XI9/XI1/XI6/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI6/MM5 N_XI9/XI1/XI6/NET44_XI9/XI1/XI6/MM5_d
+ N_X_SEL<1>_XI9/XI1/XI6/MM5_g N_XI9/XI1/XI6/NET40_XI9/XI1/XI6/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI6/MM4 N_XI9/NET5_XI9/XI1/XI6/MM4_d N_X_SEL<2>_XI9/XI1/XI6/MM4_g
+ N_XI9/XI1/XI6/NET44_XI9/XI1/XI6/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI5/MM11 N_XI9/XI1/XI5/NET030_XI9/XI1/XI5/MM11_d
+ N_WLEN_XI9/XI1/XI5/MM11_g N_VSS_XI9/XI1/XI5/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI5/MM6 N_XI9/XI1/XI5/NET40_XI9/XI1/XI5/MM6_d
+ N_X_SEL<0>_XI9/XI1/XI5/MM6_g N_XI9/XI1/XI5/NET030_XI9/XI1/XI5/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI5/MM5 N_XI9/XI1/XI5/NET44_XI9/XI1/XI5/MM5_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI5/MM5_g N_XI9/XI1/XI5/NET40_XI9/XI1/XI5/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI5/MM4 N_XI9/NET6_XI9/XI1/XI5/MM4_d N_X_SEL<2>_XI9/XI1/XI5/MM4_g
+ N_XI9/XI1/XI5/NET44_XI9/XI1/XI5/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI4/MM11 N_XI9/XI1/XI4/NET030_XI9/XI1/XI4/MM11_d
+ N_WLEN_XI9/XI1/XI4/MM11_g N_VSS_XI9/XI1/XI4/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI4/MM6 N_XI9/XI1/XI4/NET40_XI9/XI1/XI4/MM6_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI4/MM6_g N_XI9/XI1/XI4/NET030_XI9/XI1/XI4/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI4/MM5 N_XI9/XI1/XI4/NET44_XI9/XI1/XI4/MM5_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI4/MM5_g N_XI9/XI1/XI4/NET40_XI9/XI1/XI4/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI4/MM4 N_XI9/NET7_XI9/XI1/XI4/MM4_d N_X_SEL<2>_XI9/XI1/XI4/MM4_g
+ N_XI9/XI1/XI4/NET44_XI9/XI1/XI4/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI3/MM11 N_XI9/XI1/XI3/NET030_XI9/XI1/XI3/MM11_d
+ N_WLEN_XI9/XI1/XI3/MM11_g N_VSS_XI9/XI1/XI3/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI3/MM6 N_XI9/XI1/XI3/NET40_XI9/XI1/XI3/MM6_d
+ N_X_SEL<0>_XI9/XI1/XI3/MM6_g N_XI9/XI1/XI3/NET030_XI9/XI1/XI3/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI3/MM5 N_XI9/XI1/XI3/NET44_XI9/XI1/XI3/MM5_d
+ N_X_SEL<1>_XI9/XI1/XI3/MM5_g N_XI9/XI1/XI3/NET40_XI9/XI1/XI3/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI3/MM4 N_XI9/NET8_XI9/XI1/XI3/MM4_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI3/MM4_g N_XI9/XI1/XI3/NET44_XI9/XI1/XI3/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI2/MM11 N_XI9/XI1/XI2/NET030_XI9/XI1/XI2/MM11_d
+ N_WLEN_XI9/XI1/XI2/MM11_g N_VSS_XI9/XI1/XI2/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI2/MM6 N_XI9/XI1/XI2/NET40_XI9/XI1/XI2/MM6_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI2/MM6_g N_XI9/XI1/XI2/NET030_XI9/XI1/XI2/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI2/MM5 N_XI9/XI1/XI2/NET44_XI9/XI1/XI2/MM5_d
+ N_X_SEL<1>_XI9/XI1/XI2/MM5_g N_XI9/XI1/XI2/NET40_XI9/XI1/XI2/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI2/MM4 N_XI9/NET9_XI9/XI1/XI2/MM4_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI2/MM4_g N_XI9/XI1/XI2/NET44_XI9/XI1/XI2/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI1/MM11 N_XI9/XI1/XI1/NET030_XI9/XI1/XI1/MM11_d
+ N_WLEN_XI9/XI1/XI1/MM11_g N_VSS_XI9/XI1/XI1/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI1/MM6 N_XI9/XI1/XI1/NET40_XI9/XI1/XI1/MM6_d
+ N_X_SEL<0>_XI9/XI1/XI1/MM6_g N_XI9/XI1/XI1/NET030_XI9/XI1/XI1/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI1/MM5 N_XI9/XI1/XI1/NET44_XI9/XI1/XI1/MM5_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI1/MM5_g N_XI9/XI1/XI1/NET40_XI9/XI1/XI1/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI1/MM4 N_XI9/NET10_XI9/XI1/XI1/MM4_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI1/MM4_g N_XI9/XI1/XI1/NET44_XI9/XI1/XI1/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI0/MM11 N_XI9/XI1/XI0/NET030_XI9/XI1/XI0/MM11_d
+ N_WLEN_XI9/XI1/XI0/MM11_g N_VSS_XI9/XI1/XI0/MM11_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI1/XI0/MM6 N_XI9/XI1/XI0/NET40_XI9/XI1/XI0/MM6_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI0/MM6_g N_XI9/XI1/XI0/NET030_XI9/XI1/XI0/MM6_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI0/MM5 N_XI9/XI1/XI0/NET44_XI9/XI1/XI0/MM5_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI0/MM5_g N_XI9/XI1/XI0/NET40_XI9/XI1/XI0/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI1/XI0/MM4 N_XI9/NET11_XI9/XI1/XI0/MM4_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI0/MM4_g N_XI9/XI1/XI0/NET44_XI9/XI1/XI0/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI136/MM4 N_WL<63>_XI9/XI136/MM4_d N_XI9/NET4_XI9/XI136/MM4_g
+ N_VSS_XI9/XI136/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI135/MM4 N_WL<62>_XI9/XI135/MM4_d N_XI9/NET5_XI9/XI135/MM4_g
+ N_VSS_XI9/XI135/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI137/MM4 N_WL<61>_XI9/XI137/MM4_d N_XI9/NET6_XI9/XI137/MM4_g
+ N_VSS_XI9/XI137/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI138/MM4 N_WL<60>_XI9/XI138/MM4_d N_XI9/NET7_XI9/XI138/MM4_g
+ N_VSS_XI9/XI138/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI133/MM4 N_WL<59>_XI9/XI133/MM4_d N_XI9/NET8_XI9/XI133/MM4_g
+ N_VSS_XI9/XI133/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI134/MM4 N_WL<58>_XI9/XI134/MM4_d N_XI9/NET9_XI9/XI134/MM4_g
+ N_VSS_XI9/XI134/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI132/MM4 N_WL<57>_XI9/XI132/MM4_d N_XI9/NET10_XI9/XI132/MM4_g
+ N_VSS_XI9/XI132/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI131/MM4 N_WL<56>_XI9/XI131/MM4_d N_XI9/NET11_XI9/XI131/MM4_g
+ N_VSS_XI9/XI131/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI141/MM4 N_WL<55>_XI9/XI141/MM4_d N_XI9/NET4_XI9/XI141/MM4_g
+ N_VSS_XI9/XI141/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI142/MM4 N_WL<54>_XI9/XI142/MM4_d N_XI9/NET5_XI9/XI142/MM4_g
+ N_VSS_XI9/XI142/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI140/MM4 N_WL<53>_XI9/XI140/MM4_d N_XI9/NET6_XI9/XI140/MM4_g
+ N_VSS_XI9/XI140/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI139/MM4 N_WL<52>_XI9/XI139/MM4_d N_XI9/NET7_XI9/XI139/MM4_g
+ N_VSS_XI9/XI139/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI144/MM4 N_WL<51>_XI9/XI144/MM4_d N_XI9/NET8_XI9/XI144/MM4_g
+ N_VSS_XI9/XI144/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI143/MM4 N_WL<50>_XI9/XI143/MM4_d N_XI9/NET9_XI9/XI143/MM4_g
+ N_VSS_XI9/XI143/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI145/MM4 N_WL<49>_XI9/XI145/MM4_d N_XI9/NET10_XI9/XI145/MM4_g
+ N_VSS_XI9/XI145/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI146/MM4 N_WL<48>_XI9/XI146/MM4_d N_XI9/NET11_XI9/XI146/MM4_g
+ N_VSS_XI9/XI146/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI125/MM4 N_WL<47>_XI9/XI125/MM4_d N_XI9/NET4_XI9/XI125/MM4_g
+ N_VSS_XI9/XI125/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI126/MM4 N_WL<46>_XI9/XI126/MM4_d N_XI9/NET5_XI9/XI126/MM4_g
+ N_VSS_XI9/XI126/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI124/MM4 N_WL<45>_XI9/XI124/MM4_d N_XI9/NET6_XI9/XI124/MM4_g
+ N_VSS_XI9/XI124/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI123/MM4 N_WL<44>_XI9/XI123/MM4_d N_XI9/NET7_XI9/XI123/MM4_g
+ N_VSS_XI9/XI123/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI128/MM4 N_WL<43>_XI9/XI128/MM4_d N_XI9/NET8_XI9/XI128/MM4_g
+ N_VSS_XI9/XI128/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI127/MM4 N_WL<42>_XI9/XI127/MM4_d N_XI9/NET9_XI9/XI127/MM4_g
+ N_VSS_XI9/XI127/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI129/MM4 N_WL<41>_XI9/XI129/MM4_d N_XI9/NET10_XI9/XI129/MM4_g
+ N_VSS_XI9/XI129/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI130/MM4 N_WL<40>_XI9/XI130/MM4_d N_XI9/NET11_XI9/XI130/MM4_g
+ N_VSS_XI9/XI130/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI120/MM4 N_WL<39>_XI9/XI120/MM4_d N_XI9/NET4_XI9/XI120/MM4_g
+ N_VSS_XI9/XI120/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI119/MM4 N_WL<38>_XI9/XI119/MM4_d N_XI9/NET5_XI9/XI119/MM4_g
+ N_VSS_XI9/XI119/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI121/MM4 N_WL<37>_XI9/XI121/MM4_d N_XI9/NET6_XI9/XI121/MM4_g
+ N_VSS_XI9/XI121/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI122/MM4 N_WL<36>_XI9/XI122/MM4_d N_XI9/NET7_XI9/XI122/MM4_g
+ N_VSS_XI9/XI122/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI117/MM4 N_WL<35>_XI9/XI117/MM4_d N_XI9/NET8_XI9/XI117/MM4_g
+ N_VSS_XI9/XI117/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI118/MM4 N_WL<34>_XI9/XI118/MM4_d N_XI9/NET9_XI9/XI118/MM4_g
+ N_VSS_XI9/XI118/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI116/MM4 N_WL<33>_XI9/XI116/MM4_d N_XI9/NET10_XI9/XI116/MM4_g
+ N_VSS_XI9/XI116/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI115/MM4 N_WL<32>_XI9/XI115/MM4_d N_XI9/NET11_XI9/XI115/MM4_g
+ N_VSS_XI9/XI115/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI104/MM4 N_WL<31>_XI9/XI104/MM4_d N_XI9/NET4_XI9/XI104/MM4_g
+ N_VSS_XI9/XI104/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI103/MM4 N_WL<30>_XI9/XI103/MM4_d N_XI9/NET5_XI9/XI103/MM4_g
+ N_VSS_XI9/XI103/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI105/MM4 N_WL<29>_XI9/XI105/MM4_d N_XI9/NET6_XI9/XI105/MM4_g
+ N_VSS_XI9/XI105/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI106/MM4 N_WL<28>_XI9/XI106/MM4_d N_XI9/NET7_XI9/XI106/MM4_g
+ N_VSS_XI9/XI106/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI101/MM4 N_WL<27>_XI9/XI101/MM4_d N_XI9/NET8_XI9/XI101/MM4_g
+ N_VSS_XI9/XI101/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI102/MM4 N_WL<26>_XI9/XI102/MM4_d N_XI9/NET9_XI9/XI102/MM4_g
+ N_VSS_XI9/XI102/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI100/MM4 N_WL<25>_XI9/XI100/MM4_d N_XI9/NET10_XI9/XI100/MM4_g
+ N_VSS_XI9/XI100/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI99/MM4 N_WL<24>_XI9/XI99/MM4_d N_XI9/NET11_XI9/XI99/MM4_g
+ N_VSS_XI9/XI99/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI109/MM4 N_WL<23>_XI9/XI109/MM4_d N_XI9/NET4_XI9/XI109/MM4_g
+ N_VSS_XI9/XI109/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI110/MM4 N_WL<22>_XI9/XI110/MM4_d N_XI9/NET5_XI9/XI110/MM4_g
+ N_VSS_XI9/XI110/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI108/MM4 N_WL<21>_XI9/XI108/MM4_d N_XI9/NET6_XI9/XI108/MM4_g
+ N_VSS_XI9/XI108/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI107/MM4 N_WL<20>_XI9/XI107/MM4_d N_XI9/NET7_XI9/XI107/MM4_g
+ N_VSS_XI9/XI107/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI112/MM4 N_WL<19>_XI9/XI112/MM4_d N_XI9/NET8_XI9/XI112/MM4_g
+ N_VSS_XI9/XI112/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI111/MM4 N_WL<18>_XI9/XI111/MM4_d N_XI9/NET9_XI9/XI111/MM4_g
+ N_VSS_XI9/XI111/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI113/MM4 N_WL<17>_XI9/XI113/MM4_d N_XI9/NET10_XI9/XI113/MM4_g
+ N_VSS_XI9/XI113/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI114/MM4 N_WL<16>_XI9/XI114/MM4_d N_XI9/NET11_XI9/XI114/MM4_g
+ N_VSS_XI9/XI114/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI93/MM4 N_WL<15>_XI9/XI93/MM4_d N_XI9/NET4_XI9/XI93/MM4_g
+ N_VSS_XI9/XI93/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI94/MM4 N_WL<14>_XI9/XI94/MM4_d N_XI9/NET5_XI9/XI94/MM4_g
+ N_VSS_XI9/XI94/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI92/MM4 N_WL<13>_XI9/XI92/MM4_d N_XI9/NET6_XI9/XI92/MM4_g
+ N_VSS_XI9/XI92/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI91/MM4 N_WL<12>_XI9/XI91/MM4_d N_XI9/NET7_XI9/XI91/MM4_g
+ N_VSS_XI9/XI91/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI96/MM4 N_WL<11>_XI9/XI96/MM4_d N_XI9/NET8_XI9/XI96/MM4_g
+ N_VSS_XI9/XI96/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI95/MM4 N_WL<10>_XI9/XI95/MM4_d N_XI9/NET9_XI9/XI95/MM4_g
+ N_VSS_XI9/XI95/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI97/MM4 N_WL<9>_XI9/XI97/MM4_d N_XI9/NET10_XI9/XI97/MM4_g
+ N_VSS_XI9/XI97/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI98/MM4 N_WL<8>_XI9/XI98/MM4_d N_XI9/NET11_XI9/XI98/MM4_g
+ N_VSS_XI9/XI98/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI88/MM4 N_WL<7>_XI9/XI88/MM4_d N_XI9/NET4_XI9/XI88/MM4_g
+ N_VSS_XI9/XI88/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI87/MM4 N_WL<6>_XI9/XI87/MM4_d N_XI9/NET5_XI9/XI87/MM4_g
+ N_VSS_XI9/XI87/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI89/MM4 N_WL<5>_XI9/XI89/MM4_d N_XI9/NET6_XI9/XI89/MM4_g
+ N_VSS_XI9/XI89/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI90/MM4 N_WL<4>_XI9/XI90/MM4_d N_XI9/NET7_XI9/XI90/MM4_g
+ N_VSS_XI9/XI90/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI85/MM4 N_WL<3>_XI9/XI85/MM4_d N_XI9/NET8_XI9/XI85/MM4_g
+ N_VSS_XI9/XI85/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI86/MM4 N_WL<2>_XI9/XI86/MM4_d N_XI9/NET9_XI9/XI86/MM4_g
+ N_VSS_XI9/XI86/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI84/MM4 N_WL<1>_XI9/XI84/MM4_d N_XI9/NET10_XI9/XI84/MM4_g
+ N_VSS_XI9/XI84/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI2/MM4 N_WL<0>_XI9/XI2/MM4_d N_XI9/NET11_XI9/XI2/MM4_g N_VSS_XI9/XI2/MM4_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI9/XI136/MM5 N_WL<63>_XI9/XI136/MM5_d N_XI9/NET17_XI9/XI136/MM5_g
+ N_VSS_XI9/XI136/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI135/MM5 N_WL<62>_XI9/XI135/MM5_d N_XI9/NET17_XI9/XI135/MM5_g
+ N_VSS_XI9/XI135/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI137/MM5 N_WL<61>_XI9/XI137/MM5_d N_XI9/NET17_XI9/XI137/MM5_g
+ N_VSS_XI9/XI137/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI138/MM5 N_WL<60>_XI9/XI138/MM5_d N_XI9/NET17_XI9/XI138/MM5_g
+ N_VSS_XI9/XI138/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI133/MM5 N_WL<59>_XI9/XI133/MM5_d N_XI9/NET17_XI9/XI133/MM5_g
+ N_VSS_XI9/XI133/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI134/MM5 N_WL<58>_XI9/XI134/MM5_d N_XI9/NET17_XI9/XI134/MM5_g
+ N_VSS_XI9/XI134/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI132/MM5 N_WL<57>_XI9/XI132/MM5_d N_XI9/NET17_XI9/XI132/MM5_g
+ N_VSS_XI9/XI132/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI131/MM5 N_WL<56>_XI9/XI131/MM5_d N_XI9/NET17_XI9/XI131/MM5_g
+ N_VSS_XI9/XI131/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI141/MM5 N_WL<55>_XI9/XI141/MM5_d N_XI9/NET18_XI9/XI141/MM5_g
+ N_VSS_XI9/XI141/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI142/MM5 N_WL<54>_XI9/XI142/MM5_d N_XI9/NET18_XI9/XI142/MM5_g
+ N_VSS_XI9/XI142/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI140/MM5 N_WL<53>_XI9/XI140/MM5_d N_XI9/NET18_XI9/XI140/MM5_g
+ N_VSS_XI9/XI140/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI139/MM5 N_WL<52>_XI9/XI139/MM5_d N_XI9/NET18_XI9/XI139/MM5_g
+ N_VSS_XI9/XI139/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI144/MM5 N_WL<51>_XI9/XI144/MM5_d N_XI9/NET18_XI9/XI144/MM5_g
+ N_VSS_XI9/XI144/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI143/MM5 N_WL<50>_XI9/XI143/MM5_d N_XI9/NET18_XI9/XI143/MM5_g
+ N_VSS_XI9/XI143/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI145/MM5 N_WL<49>_XI9/XI145/MM5_d N_XI9/NET18_XI9/XI145/MM5_g
+ N_VSS_XI9/XI145/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI146/MM5 N_WL<48>_XI9/XI146/MM5_d N_XI9/NET18_XI9/XI146/MM5_g
+ N_VSS_XI9/XI146/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI125/MM5 N_WL<47>_XI9/XI125/MM5_d N_XI9/NET19_XI9/XI125/MM5_g
+ N_VSS_XI9/XI125/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI126/MM5 N_WL<46>_XI9/XI126/MM5_d N_XI9/NET19_XI9/XI126/MM5_g
+ N_VSS_XI9/XI126/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI124/MM5 N_WL<45>_XI9/XI124/MM5_d N_XI9/NET19_XI9/XI124/MM5_g
+ N_VSS_XI9/XI124/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI123/MM5 N_WL<44>_XI9/XI123/MM5_d N_XI9/NET19_XI9/XI123/MM5_g
+ N_VSS_XI9/XI123/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI128/MM5 N_WL<43>_XI9/XI128/MM5_d N_XI9/NET19_XI9/XI128/MM5_g
+ N_VSS_XI9/XI128/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI127/MM5 N_WL<42>_XI9/XI127/MM5_d N_XI9/NET19_XI9/XI127/MM5_g
+ N_VSS_XI9/XI127/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI129/MM5 N_WL<41>_XI9/XI129/MM5_d N_XI9/NET19_XI9/XI129/MM5_g
+ N_VSS_XI9/XI129/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI130/MM5 N_WL<40>_XI9/XI130/MM5_d N_XI9/NET19_XI9/XI130/MM5_g
+ N_VSS_XI9/XI130/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI120/MM5 N_WL<39>_XI9/XI120/MM5_d N_XI9/NET20_XI9/XI120/MM5_g
+ N_VSS_XI9/XI120/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI119/MM5 N_WL<38>_XI9/XI119/MM5_d N_XI9/NET20_XI9/XI119/MM5_g
+ N_VSS_XI9/XI119/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI121/MM5 N_WL<37>_XI9/XI121/MM5_d N_XI9/NET20_XI9/XI121/MM5_g
+ N_VSS_XI9/XI121/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI122/MM5 N_WL<36>_XI9/XI122/MM5_d N_XI9/NET20_XI9/XI122/MM5_g
+ N_VSS_XI9/XI122/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI117/MM5 N_WL<35>_XI9/XI117/MM5_d N_XI9/NET20_XI9/XI117/MM5_g
+ N_VSS_XI9/XI117/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI118/MM5 N_WL<34>_XI9/XI118/MM5_d N_XI9/NET20_XI9/XI118/MM5_g
+ N_VSS_XI9/XI118/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI116/MM5 N_WL<33>_XI9/XI116/MM5_d N_XI9/NET20_XI9/XI116/MM5_g
+ N_VSS_XI9/XI116/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI115/MM5 N_WL<32>_XI9/XI115/MM5_d N_XI9/NET20_XI9/XI115/MM5_g
+ N_VSS_XI9/XI115/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI104/MM5 N_WL<31>_XI9/XI104/MM5_d N_XI9/NET21_XI9/XI104/MM5_g
+ N_VSS_XI9/XI104/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI103/MM5 N_WL<30>_XI9/XI103/MM5_d N_XI9/NET21_XI9/XI103/MM5_g
+ N_VSS_XI9/XI103/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI105/MM5 N_WL<29>_XI9/XI105/MM5_d N_XI9/NET21_XI9/XI105/MM5_g
+ N_VSS_XI9/XI105/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI106/MM5 N_WL<28>_XI9/XI106/MM5_d N_XI9/NET21_XI9/XI106/MM5_g
+ N_VSS_XI9/XI106/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI101/MM5 N_WL<27>_XI9/XI101/MM5_d N_XI9/NET21_XI9/XI101/MM5_g
+ N_VSS_XI9/XI101/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI102/MM5 N_WL<26>_XI9/XI102/MM5_d N_XI9/NET21_XI9/XI102/MM5_g
+ N_VSS_XI9/XI102/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI100/MM5 N_WL<25>_XI9/XI100/MM5_d N_XI9/NET21_XI9/XI100/MM5_g
+ N_VSS_XI9/XI100/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI99/MM5 N_WL<24>_XI9/XI99/MM5_d N_XI9/NET21_XI9/XI99/MM5_g
+ N_VSS_XI9/XI99/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI109/MM5 N_WL<23>_XI9/XI109/MM5_d N_XI9/NET22_XI9/XI109/MM5_g
+ N_VSS_XI9/XI109/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI110/MM5 N_WL<22>_XI9/XI110/MM5_d N_XI9/NET22_XI9/XI110/MM5_g
+ N_VSS_XI9/XI110/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI108/MM5 N_WL<21>_XI9/XI108/MM5_d N_XI9/NET22_XI9/XI108/MM5_g
+ N_VSS_XI9/XI108/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI107/MM5 N_WL<20>_XI9/XI107/MM5_d N_XI9/NET22_XI9/XI107/MM5_g
+ N_VSS_XI9/XI107/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI112/MM5 N_WL<19>_XI9/XI112/MM5_d N_XI9/NET22_XI9/XI112/MM5_g
+ N_VSS_XI9/XI112/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI111/MM5 N_WL<18>_XI9/XI111/MM5_d N_XI9/NET22_XI9/XI111/MM5_g
+ N_VSS_XI9/XI111/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI113/MM5 N_WL<17>_XI9/XI113/MM5_d N_XI9/NET22_XI9/XI113/MM5_g
+ N_VSS_XI9/XI113/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI114/MM5 N_WL<16>_XI9/XI114/MM5_d N_XI9/NET22_XI9/XI114/MM5_g
+ N_VSS_XI9/XI114/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI93/MM5 N_WL<15>_XI9/XI93/MM5_d N_XI9/NET23_XI9/XI93/MM5_g
+ N_VSS_XI9/XI93/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI94/MM5 N_WL<14>_XI9/XI94/MM5_d N_XI9/NET23_XI9/XI94/MM5_g
+ N_VSS_XI9/XI94/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI92/MM5 N_WL<13>_XI9/XI92/MM5_d N_XI9/NET23_XI9/XI92/MM5_g
+ N_VSS_XI9/XI92/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI91/MM5 N_WL<12>_XI9/XI91/MM5_d N_XI9/NET23_XI9/XI91/MM5_g
+ N_VSS_XI9/XI91/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI96/MM5 N_WL<11>_XI9/XI96/MM5_d N_XI9/NET23_XI9/XI96/MM5_g
+ N_VSS_XI9/XI96/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI95/MM5 N_WL<10>_XI9/XI95/MM5_d N_XI9/NET23_XI9/XI95/MM5_g
+ N_VSS_XI9/XI95/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI97/MM5 N_WL<9>_XI9/XI97/MM5_d N_XI9/NET23_XI9/XI97/MM5_g
+ N_VSS_XI9/XI97/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI98/MM5 N_WL<8>_XI9/XI98/MM5_d N_XI9/NET23_XI9/XI98/MM5_g
+ N_VSS_XI9/XI98/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI88/MM5 N_WL<7>_XI9/XI88/MM5_d N_XI9/NET24_XI9/XI88/MM5_g
+ N_VSS_XI9/XI88/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI87/MM5 N_WL<6>_XI9/XI87/MM5_d N_XI9/NET24_XI9/XI87/MM5_g
+ N_VSS_XI9/XI87/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI89/MM5 N_WL<5>_XI9/XI89/MM5_d N_XI9/NET24_XI9/XI89/MM5_g
+ N_VSS_XI9/XI89/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI90/MM5 N_WL<4>_XI9/XI90/MM5_d N_XI9/NET24_XI9/XI90/MM5_g
+ N_VSS_XI9/XI90/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI85/MM5 N_WL<3>_XI9/XI85/MM5_d N_XI9/NET24_XI9/XI85/MM5_g
+ N_VSS_XI9/XI85/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI86/MM5 N_WL<2>_XI9/XI86/MM5_d N_XI9/NET24_XI9/XI86/MM5_g
+ N_VSS_XI9/XI86/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI84/MM5 N_WL<1>_XI9/XI84/MM5_d N_XI9/NET24_XI9/XI84/MM5_g
+ N_VSS_XI9/XI84/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9/XI2/MM5 N_WL<0>_XI9/XI2/MM5_d N_XI9/NET24_XI9/XI2/MM5_g N_VSS_XI9/XI2/MM5_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI10/MM2460 N_VSS_XI10/MM2460_d N_WL<63>_XI10/MM2460_g N_BL<0>_XI10/MM2460_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2418 N_VSS_XI10/MM2418_d N_WL<62>_XI10/MM2418_g XI10/NET3768
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2499 N_VSS_XI10/MM2499_d N_WL<61>_XI10/MM2499_g N_BL<0>_XI10/MM2499_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2532 N_VSS_XI10/MM2532_d N_WL<60>_XI10/MM2532_g XI10/NET5060
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2344 N_VSS_XI10/MM2344_d N_WL<59>_XI10/MM2344_g N_BL<0>_XI10/MM2344_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2376 N_VSS_XI10/MM2376_d N_WL<58>_XI10/MM2376_g XI10/NET3860
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2563 N_VSS_XI10/MM2563_d N_WL<57>_XI10/MM2563_g N_BL<0>_XI10/MM2563_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2496 N_VSS_XI10/MM2496_d N_WL<56>_XI10/MM2496_g XI10/NET5096
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2207 N_VSS_XI10/MM2207_d N_WL<55>_XI10/MM2207_g N_BL<0>_XI10/MM2207_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2240 N_VSS_XI10/MM2240_d N_WL<54>_XI10/MM2240_g XI10/NET4104
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2168 N_VSS_XI10/MM2168_d N_WL<53>_XI10/MM2168_g N_BL<0>_XI10/MM2168_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2121 N_VSS_XI10/MM2121_d N_WL<52>_XI10/MM2121_g XI10/NET3500
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2323 N_VSS_XI10/MM2323_d N_WL<51>_XI10/MM2323_g N_BL<0>_XI10/MM2323_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2277 N_VSS_XI10/MM2277_d N_WL<50>_XI10/MM2277_g XI10/NET4032
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2104 N_VSS_XI10/MM2104_d N_WL<49>_XI10/MM2104_g N_BL<0>_XI10/MM2104_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2171 N_VSS_XI10/MM2171_d N_WL<48>_XI10/MM2171_g XI10/NET4232
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2719 N_VSS_XI10/MM2719_d N_WL<47>_XI10/MM2719_g N_BL<0>_XI10/MM2719_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2752 N_VSS_XI10/MM2752_d N_WL<46>_XI10/MM2752_g XI10/NET4572
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2680 N_VSS_XI10/MM2680_d N_WL<45>_XI10/MM2680_g N_BL<0>_XI10/MM2680_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2633 N_VSS_XI10/MM2633_d N_WL<44>_XI10/MM2633_g XI10/NET4792
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2835 N_VSS_XI10/MM2835_d N_WL<43>_XI10/MM2835_g N_BL<0>_XI10/MM2835_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2789 N_VSS_XI10/MM2789_d N_WL<42>_XI10/MM2789_g XI10/NET4500
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2616 N_VSS_XI10/MM2616_d N_WL<41>_XI10/MM2616_g N_BL<0>_XI10/MM2616_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2590 N_VSS_XI10/MM2590_d N_WL<40>_XI10/MM2590_g XI10/NET4896
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2972 N_VSS_XI10/MM2972_d N_WL<39>_XI10/MM2972_g N_BL<0>_XI10/MM2972_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2925 N_VSS_XI10/MM2925_d N_WL<38>_XI10/MM2925_g XI10/NET5456
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3011 N_VSS_XI10/MM3011_d N_WL<37>_XI10/MM3011_g N_BL<0>_XI10/MM3011_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3044 N_VSS_XI10/MM3044_d N_WL<36>_XI10/MM3044_g XI10/NET5236
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2856 N_VSS_XI10/MM2856_d N_WL<35>_XI10/MM2856_g N_BL<0>_XI10/MM2856_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2888 N_VSS_XI10/MM2888_d N_WL<34>_XI10/MM2888_g XI10/NET4328
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3075 N_VSS_XI10/MM3075_d N_WL<33>_XI10/MM3075_g N_BL<0>_XI10/MM3075_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3085 N_VSS_XI10/MM3085_d N_WL<32>_XI10/MM3085_g XI10/NET5484
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1695 N_VSS_XI10/MM1695_d N_WL<31>_XI10/MM1695_g N_BL<0>_XI10/MM1695_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1728 N_VSS_XI10/MM1728_d N_WL<30>_XI10/MM1728_g XI10/NET2136
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1656 N_VSS_XI10/MM1656_d N_WL<29>_XI10/MM1656_g N_BL<0>_XI10/MM1656_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1609 N_VSS_XI10/MM1609_d N_WL<28>_XI10/MM1609_g XI10/NET2356
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1811 N_VSS_XI10/MM1811_d N_WL<27>_XI10/MM1811_g N_BL<0>_XI10/MM1811_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1765 N_VSS_XI10/MM1765_d N_WL<26>_XI10/MM1765_g XI10/NET2064
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1592 N_VSS_XI10/MM1592_d N_WL<25>_XI10/MM1592_g N_BL<0>_XI10/MM1592_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1566 N_VSS_XI10/MM1566_d N_WL<24>_XI10/MM1566_g XI10/NET2460
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1948 N_VSS_XI10/MM1948_d N_WL<23>_XI10/MM1948_g N_BL<0>_XI10/MM1948_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1901 N_VSS_XI10/MM1901_d N_WL<22>_XI10/MM1901_g XI10/NET2844
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1987 N_VSS_XI10/MM1987_d N_WL<21>_XI10/MM1987_g N_BL<0>_XI10/MM1987_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2020 N_VSS_XI10/MM2020_d N_WL<20>_XI10/MM2020_g XI10/NET02641
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1832 N_VSS_XI10/MM1832_d N_WL<19>_XI10/MM1832_g N_BL<0>_XI10/MM1832_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1864 N_VSS_XI10/MM1864_d N_WL<18>_XI10/MM1864_g XI10/NET2916
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2051 N_VSS_XI10/MM2051_d N_WL<17>_XI10/MM2051_g N_BL<0>_XI10/MM2051_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1900 N_VSS_XI10/MM1900_d N_WL<16>_XI10/MM1900_g XI10/NET2848
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1436 N_VSS_XI10/MM1436_d N_WL<15>_XI10/MM1436_g N_BL<0>_XI10/MM1436_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1403 N_VSS_XI10/MM1403_d N_WL<14>_XI10/MM1403_g XI10/NET5632
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1475 N_VSS_XI10/MM1475_d N_WL<13>_XI10/MM1475_g N_BL<0>_XI10/MM1475_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1508 N_VSS_XI10/MM1508_d N_WL<12>_XI10/MM1508_g XI10/NET1872
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1320 N_VSS_XI10/MM1320_d N_WL<11>_XI10/MM1320_g N_BL<0>_XI10/MM1320_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1366 N_VSS_XI10/MM1366_d N_WL<10>_XI10/MM1366_g XI10/NET5560
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1539 N_VSS_XI10/MM1539_d N_WL<9>_XI10/MM1539_g N_BL<0>_XI10/MM1539_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1472 N_VSS_XI10/MM1472_d N_WL<8>_XI10/MM1472_g XI10/NET5764
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1228 N_VSS_XI10/MM1228_d N_WL<7>_XI10/MM1228_g N_BL<0>_XI10/MM1228_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1196 N_VSS_XI10/MM1196_d N_WL<6>_XI10/MM1196_g XI10/NET3088
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1263 N_VSS_XI10/MM1263_d N_WL<5>_XI10/MM1263_g N_BL<0>_XI10/MM1263_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1309 N_VSS_XI10/MM1309_d N_WL<4>_XI10/MM1309_g XI10/NET3308
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1135 N_VSS_XI10/MM1135_d N_WL<3>_XI10/MM1135_g N_BL<0>_XI10/MM1135_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1181 N_VSS_XI10/MM1181_d N_WL<2>_XI10/MM1181_g XI10/NET1992
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1116 N_VSS_XI10/MM1116_d N_WL<1>_XI10/MM1116_g N_BL<0>_XI10/MM1116_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM0 N_VSS_XI10/MM0_d N_WL<0>_XI10/MM0_g XI10/NET5804 N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI16/XI21/XI1/MM10 N_XI16/XI21/NET40_XI16/XI21/XI1/MM10_d
+ N_YOUT<1>_XI16/XI21/XI1/MM10_g N_VSS_XI16/XI21/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI22/XI1/MM10 N_XI16/XI22/NET40_XI16/XI22/XI1/MM10_d
+ N_YOUT<0>_XI16/XI22/XI1/MM10_g N_VSS_XI16/XI22/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI21/MM1 N_BL<1>_XI16/XI21/MM1_d N_XI16/XI21/NET40_XI16/XI21/MM1_g
+ N_DL<0>_XI16/XI21/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI22/MM1 N_BL<0>_XI16/XI22/MM1_d N_XI16/XI22/NET40_XI16/XI22/MM1_g
+ N_DL<0>_XI16/XI22/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2447 N_VSS_XI10/MM2447_d N_WL<63>_XI10/MM2447_g XI10/NET3720
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2414 N_VSS_XI10/MM2414_d N_WL<62>_XI10/MM2414_g N_BL<1>_XI10/MM2414_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2497 N_VSS_XI10/MM2497_d N_WL<61>_XI10/MM2497_g XI10/NET5092
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2545 N_VSS_XI10/MM2545_d N_WL<60>_XI10/MM2545_g N_BL<1>_XI10/MM2545_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2564 N_VSS_XI10/MM2564_d N_WL<59>_XI10/MM2564_g XI10/NET4936
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2389 N_VSS_XI10/MM2389_d N_WL<58>_XI10/MM2389_g N_BL<1>_XI10/MM2389_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2556 N_VSS_XI10/MM2556_d N_WL<57>_XI10/MM2556_g XI10/NET4968
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2588 N_VSS_XI10/MM2588_d N_WL<56>_XI10/MM2588_g N_BL<1>_XI10/MM2588_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2195 N_VSS_XI10/MM2195_d N_WL<55>_XI10/MM2195_g XI10/NET4172
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2253 N_VSS_XI10/MM2253_d N_WL<54>_XI10/MM2253_g N_BL<1>_XI10/MM2253_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2154 N_VSS_XI10/MM2154_d N_WL<53>_XI10/MM2154_g XI10/NET4260
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2122 N_VSS_XI10/MM2122_d N_WL<52>_XI10/MM2122_g N_BL<1>_XI10/MM2122_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2310 N_VSS_XI10/MM2310_d N_WL<51>_XI10/MM2310_g XI10/NET3968
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2278 N_VSS_XI10/MM2278_d N_WL<50>_XI10/MM2278_g N_BL<1>_XI10/MM2278_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2231 N_VSS_XI10/MM2231_d N_WL<49>_XI10/MM2231_g XI10/NET4112
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2079 N_VSS_XI10/MM2079_d N_WL<48>_XI10/MM2079_g N_BL<1>_XI10/MM2079_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2707 N_VSS_XI10/MM2707_d N_WL<47>_XI10/MM2707_g XI10/NET4640
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2765 N_VSS_XI10/MM2765_d N_WL<46>_XI10/MM2765_g N_BL<1>_XI10/MM2765_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2666 N_VSS_XI10/MM2666_d N_WL<45>_XI10/MM2666_g XI10/NET4728
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2634 N_VSS_XI10/MM2634_d N_WL<44>_XI10/MM2634_g N_BL<1>_XI10/MM2634_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2609 N_VSS_XI10/MM2609_d N_WL<43>_XI10/MM2609_g XI10/NET4876
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2790 N_VSS_XI10/MM2790_d N_WL<42>_XI10/MM2790_g N_BL<1>_XI10/MM2790_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2593 N_VSS_XI10/MM2593_d N_WL<41>_XI10/MM2593_g XI10/NET4888
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2591 N_VSS_XI10/MM2591_d N_WL<40>_XI10/MM2591_g N_BL<1>_XI10/MM2591_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2959 N_VSS_XI10/MM2959_d N_WL<39>_XI10/MM2959_g XI10/NET5388
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2926 N_VSS_XI10/MM2926_d N_WL<38>_XI10/MM2926_g N_BL<1>_XI10/MM2926_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2995 N_VSS_XI10/MM2995_d N_WL<37>_XI10/MM2995_g XI10/NET5320
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3057 N_VSS_XI10/MM3057_d N_WL<36>_XI10/MM3057_g N_BL<1>_XI10/MM3057_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3082 N_VSS_XI10/MM3082_d N_WL<35>_XI10/MM3082_g XI10/NET5488
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2901 N_VSS_XI10/MM2901_d N_WL<34>_XI10/MM2901_g N_BL<1>_XI10/MM2901_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3098 N_VSS_XI10/MM3098_d N_WL<33>_XI10/MM3098_g XI10/NET5476
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3100 N_VSS_XI10/MM3100_d N_WL<32>_XI10/MM3100_g N_BL<1>_XI10/MM3100_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1683 N_VSS_XI10/MM1683_d N_WL<31>_XI10/MM1683_g XI10/NET2204
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1741 N_VSS_XI10/MM1741_d N_WL<30>_XI10/MM1741_g N_BL<1>_XI10/MM1741_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1642 N_VSS_XI10/MM1642_d N_WL<29>_XI10/MM1642_g XI10/NET2292
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1610 N_VSS_XI10/MM1610_d N_WL<28>_XI10/MM1610_g N_BL<1>_XI10/MM1610_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1810 N_VSS_XI10/MM1810_d N_WL<27>_XI10/MM1810_g XI10/NET3016
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1766 N_VSS_XI10/MM1766_d N_WL<26>_XI10/MM1766_g N_BL<1>_XI10/MM1766_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1569 N_VSS_XI10/MM1569_d N_WL<25>_XI10/MM1569_g XI10/NET2452
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1567 N_VSS_XI10/MM1567_d N_WL<24>_XI10/MM1567_g N_BL<1>_XI10/MM1567_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1935 N_VSS_XI10/MM1935_d N_WL<23>_XI10/MM1935_g XI10/NET2776
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1902 N_VSS_XI10/MM1902_d N_WL<22>_XI10/MM1902_g N_BL<1>_XI10/MM1902_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1971 N_VSS_XI10/MM1971_d N_WL<21>_XI10/MM1971_g XI10/NET2708
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2033 N_VSS_XI10/MM2033_d N_WL<20>_XI10/MM2033_g N_BL<1>_XI10/MM2033_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1825 N_VSS_XI10/MM1825_d N_WL<19>_XI10/MM1825_g XI10/NET2964
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1877 N_VSS_XI10/MM1877_d N_WL<18>_XI10/MM1877_g N_BL<1>_XI10/MM1877_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1890 N_VSS_XI10/MM1890_d N_WL<17>_XI10/MM1890_g XI10/NET2856
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2076 N_VSS_XI10/MM2076_d N_WL<16>_XI10/MM2076_g N_BL<1>_XI10/MM2076_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1448 N_VSS_XI10/MM1448_d N_WL<15>_XI10/MM1448_g XI10/NET5700
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1390 N_VSS_XI10/MM1390_d N_WL<14>_XI10/MM1390_g N_BL<1>_XI10/MM1390_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1489 N_VSS_XI10/MM1489_d N_WL<13>_XI10/MM1489_g XI10/NET5792
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1521 N_VSS_XI10/MM1521_d N_WL<12>_XI10/MM1521_g N_BL<1>_XI10/MM1521_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1333 N_VSS_XI10/MM1333_d N_WL<11>_XI10/MM1333_g XI10/NET5496
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1365 N_VSS_XI10/MM1365_d N_WL<10>_XI10/MM1365_g N_BL<1>_XI10/MM1365_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1412 N_VSS_XI10/MM1412_d N_WL<9>_XI10/MM1412_g XI10/NET5640
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1564 N_VSS_XI10/MM1564_d N_WL<8>_XI10/MM1564_g N_BL<1>_XI10/MM1564_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1240 N_VSS_XI10/MM1240_d N_WL<7>_XI10/MM1240_g XI10/NET3156
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1183 N_VSS_XI10/MM1183_d N_WL<6>_XI10/MM1183_g N_BL<1>_XI10/MM1183_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1276 N_VSS_XI10/MM1276_d N_WL<5>_XI10/MM1276_g XI10/NET3244
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1308 N_VSS_XI10/MM1308_d N_WL<4>_XI10/MM1308_g N_BL<1>_XI10/MM1308_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1124 N_VSS_XI10/MM1124_d N_WL<3>_XI10/MM1124_g XI10/NET3436
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1180 N_VSS_XI10/MM1180_d N_WL<2>_XI10/MM1180_g N_BL<1>_XI10/MM1180_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1102 N_VSS_XI10/MM1102_d N_WL<1>_XI10/MM1102_g XI10/NET5796
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1 N_VSS_XI10/MM1_d N_WL<0>_XI10/MM1_g N_BL<1>_XI10/MM1_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2461 N_VSS_XI10/MM2461_d N_WL<63>_XI10/MM2461_g N_BL<2>_XI10/MM2461_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2427 N_VSS_XI10/MM2427_d N_WL<62>_XI10/MM2427_g XI10/NET3732
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2498 N_VSS_XI10/MM2498_d N_WL<61>_XI10/MM2498_g N_BL<2>_XI10/MM2498_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2533 N_VSS_XI10/MM2533_d N_WL<60>_XI10/MM2533_g XI10/NET5056
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2343 N_VSS_XI10/MM2343_d N_WL<59>_XI10/MM2343_g N_BL<2>_XI10/MM2343_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2377 N_VSS_XI10/MM2377_d N_WL<58>_XI10/MM2377_g XI10/NET3856
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2562 N_VSS_XI10/MM2562_d N_WL<57>_XI10/MM2562_g N_BL<2>_XI10/MM2562_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2547 N_VSS_XI10/MM2547_d N_WL<56>_XI10/MM2547_g XI10/NET5000
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2206 N_VSS_XI10/MM2206_d N_WL<55>_XI10/MM2206_g N_BL<2>_XI10/MM2206_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2241 N_VSS_XI10/MM2241_d N_WL<54>_XI10/MM2241_g XI10/NET4100
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2169 N_VSS_XI10/MM2169_d N_WL<53>_XI10/MM2169_g N_BL<2>_XI10/MM2169_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2123 N_VSS_XI10/MM2123_d N_WL<52>_XI10/MM2123_g XI10/NET3492
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2324 N_VSS_XI10/MM2324_d N_WL<51>_XI10/MM2324_g N_BL<2>_XI10/MM2324_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2279 N_VSS_XI10/MM2279_d N_WL<50>_XI10/MM2279_g XI10/NET4024
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2105 N_VSS_XI10/MM2105_d N_WL<49>_XI10/MM2105_g N_BL<2>_XI10/MM2105_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2182 N_VSS_XI10/MM2182_d N_WL<48>_XI10/MM2182_g XI10/NET4192
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2718 N_VSS_XI10/MM2718_d N_WL<47>_XI10/MM2718_g N_BL<2>_XI10/MM2718_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2753 N_VSS_XI10/MM2753_d N_WL<46>_XI10/MM2753_g XI10/NET4568
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2681 N_VSS_XI10/MM2681_d N_WL<45>_XI10/MM2681_g N_BL<2>_XI10/MM2681_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2635 N_VSS_XI10/MM2635_d N_WL<44>_XI10/MM2635_g XI10/NET4784
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2836 N_VSS_XI10/MM2836_d N_WL<43>_XI10/MM2836_g N_BL<2>_XI10/MM2836_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2791 N_VSS_XI10/MM2791_d N_WL<42>_XI10/MM2791_g XI10/NET4492
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2617 N_VSS_XI10/MM2617_d N_WL<41>_XI10/MM2617_g N_BL<2>_XI10/MM2617_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2606 N_VSS_XI10/MM2606_d N_WL<40>_XI10/MM2606_g XI10/NET4880
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2973 N_VSS_XI10/MM2973_d N_WL<39>_XI10/MM2973_g N_BL<2>_XI10/MM2973_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2927 N_VSS_XI10/MM2927_d N_WL<38>_XI10/MM2927_g XI10/NET5448
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3010 N_VSS_XI10/MM3010_d N_WL<37>_XI10/MM3010_g N_BL<2>_XI10/MM3010_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3045 N_VSS_XI10/MM3045_d N_WL<36>_XI10/MM3045_g XI10/NET5232
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2855 N_VSS_XI10/MM2855_d N_WL<35>_XI10/MM2855_g N_BL<2>_XI10/MM2855_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2889 N_VSS_XI10/MM2889_d N_WL<34>_XI10/MM2889_g XI10/NET4324
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3074 N_VSS_XI10/MM3074_d N_WL<33>_XI10/MM3074_g N_BL<2>_XI10/MM3074_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3101 N_VSS_XI10/MM3101_d N_WL<32>_XI10/MM3101_g XI10/NET5468
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1694 N_VSS_XI10/MM1694_d N_WL<31>_XI10/MM1694_g N_BL<2>_XI10/MM1694_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1729 N_VSS_XI10/MM1729_d N_WL<30>_XI10/MM1729_g XI10/NET2132
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1657 N_VSS_XI10/MM1657_d N_WL<29>_XI10/MM1657_g N_BL<2>_XI10/MM1657_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1611 N_VSS_XI10/MM1611_d N_WL<28>_XI10/MM1611_g XI10/NET2348
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1812 N_VSS_XI10/MM1812_d N_WL<27>_XI10/MM1812_g N_BL<2>_XI10/MM1812_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1767 N_VSS_XI10/MM1767_d N_WL<26>_XI10/MM1767_g XI10/NET2056
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1593 N_VSS_XI10/MM1593_d N_WL<25>_XI10/MM1593_g N_BL<2>_XI10/MM1593_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1582 N_VSS_XI10/MM1582_d N_WL<24>_XI10/MM1582_g XI10/NET2444
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1949 N_VSS_XI10/MM1949_d N_WL<23>_XI10/MM1949_g N_BL<2>_XI10/MM1949_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1903 N_VSS_XI10/MM1903_d N_WL<22>_XI10/MM1903_g XI10/NET2836
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1986 N_VSS_XI10/MM1986_d N_WL<21>_XI10/MM1986_g N_BL<2>_XI10/MM1986_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2021 N_VSS_XI10/MM2021_d N_WL<20>_XI10/MM2021_g XI10/NET02644
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1831 N_VSS_XI10/MM1831_d N_WL<19>_XI10/MM1831_g N_BL<2>_XI10/MM1831_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1865 N_VSS_XI10/MM1865_d N_WL<18>_XI10/MM1865_g XI10/NET2912
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2050 N_VSS_XI10/MM2050_d N_WL<17>_XI10/MM2050_g N_BL<2>_XI10/MM2050_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1973 N_VSS_XI10/MM1973_d N_WL<16>_XI10/MM1973_g XI10/NET2700
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1437 N_VSS_XI10/MM1437_d N_WL<15>_XI10/MM1437_g N_BL<2>_XI10/MM1437_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1402 N_VSS_XI10/MM1402_d N_WL<14>_XI10/MM1402_g XI10/NET5628
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1474 N_VSS_XI10/MM1474_d N_WL<13>_XI10/MM1474_g N_BL<2>_XI10/MM1474_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1509 N_VSS_XI10/MM1509_d N_WL<12>_XI10/MM1509_g XI10/NET1868
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1319 N_VSS_XI10/MM1319_d N_WL<11>_XI10/MM1319_g N_BL<2>_XI10/MM1319_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1364 N_VSS_XI10/MM1364_d N_WL<10>_XI10/MM1364_g XI10/NET5552
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1538 N_VSS_XI10/MM1538_d N_WL<9>_XI10/MM1538_g N_BL<2>_XI10/MM1538_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1461 N_VSS_XI10/MM1461_d N_WL<8>_XI10/MM1461_g XI10/NET5724
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1229 N_VSS_XI10/MM1229_d N_WL<7>_XI10/MM1229_g N_BL<2>_XI10/MM1229_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1195 N_VSS_XI10/MM1195_d N_WL<6>_XI10/MM1195_g XI10/NET3084
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1262 N_VSS_XI10/MM1262_d N_WL<5>_XI10/MM1262_g N_BL<2>_XI10/MM1262_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1307 N_VSS_XI10/MM1307_d N_WL<4>_XI10/MM1307_g XI10/NET3300
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1134 N_VSS_XI10/MM1134_d N_WL<3>_XI10/MM1134_g N_BL<2>_XI10/MM1134_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1179 N_VSS_XI10/MM1179_d N_WL<2>_XI10/MM1179_g XI10/NET1984
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1115 N_VSS_XI10/MM1115_d N_WL<1>_XI10/MM1115_g N_BL<2>_XI10/MM1115_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1056 N_VSS_XI10/MM1056_d N_WL<0>_XI10/MM1056_g XI10/NET4264
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI16/XI19/XI1/MM10 N_XI16/XI19/NET40_XI16/XI19/XI1/MM10_d
+ N_YOUT<3>_XI16/XI19/XI1/MM10_g N_VSS_XI16/XI19/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI20/XI1/MM10 N_XI16/XI20/NET40_XI16/XI20/XI1/MM10_d
+ N_YOUT<2>_XI16/XI20/XI1/MM10_g N_VSS_XI16/XI20/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI19/MM1 N_BL<3>_XI16/XI19/MM1_d N_XI16/XI19/NET40_XI16/XI19/MM1_g
+ N_DL<0>_XI16/XI19/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI20/MM1 N_BL<2>_XI16/XI20/MM1_d N_XI16/XI20/NET40_XI16/XI20/MM1_g
+ N_DL<0>_XI16/XI20/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2459 N_VSS_XI10/MM2459_d N_WL<63>_XI10/MM2459_g XI10/NET3712
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2416 N_VSS_XI10/MM2416_d N_WL<62>_XI10/MM2416_g N_BL<3>_XI10/MM2416_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2500 N_VSS_XI10/MM2500_d N_WL<61>_XI10/MM2500_g XI10/NET5080
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2543 N_VSS_XI10/MM2543_d N_WL<60>_XI10/MM2543_g N_BL<3>_XI10/MM2543_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2570 N_VSS_XI10/MM2570_d N_WL<59>_XI10/MM2570_g XI10/NET4920
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2387 N_VSS_XI10/MM2387_d N_WL<58>_XI10/MM2387_g N_BL<3>_XI10/MM2387_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2557 N_VSS_XI10/MM2557_d N_WL<57>_XI10/MM2557_g XI10/NET4964
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2568 N_VSS_XI10/MM2568_d N_WL<56>_XI10/MM2568_g N_BL<3>_XI10/MM2568_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2196 N_VSS_XI10/MM2196_d N_WL<55>_XI10/MM2196_g XI10/NET4168
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2251 N_VSS_XI10/MM2251_d N_WL<54>_XI10/MM2251_g N_BL<3>_XI10/MM2251_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2167 N_VSS_XI10/MM2167_d N_WL<53>_XI10/MM2167_g XI10/NET4248
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2124 N_VSS_XI10/MM2124_d N_WL<52>_XI10/MM2124_g N_BL<3>_XI10/MM2124_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2322 N_VSS_XI10/MM2322_d N_WL<51>_XI10/MM2322_g XI10/NET3960
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2280 N_VSS_XI10/MM2280_d N_WL<50>_XI10/MM2280_g N_BL<3>_XI10/MM2280_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2265 N_VSS_XI10/MM2265_d N_WL<49>_XI10/MM2265_g XI10/NET4036
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2099 N_VSS_XI10/MM2099_d N_WL<48>_XI10/MM2099_g N_BL<3>_XI10/MM2099_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2708 N_VSS_XI10/MM2708_d N_WL<47>_XI10/MM2708_g XI10/NET4636
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2763 N_VSS_XI10/MM2763_d N_WL<46>_XI10/MM2763_g N_BL<3>_XI10/MM2763_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2679 N_VSS_XI10/MM2679_d N_WL<45>_XI10/MM2679_g XI10/NET4716
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2636 N_VSS_XI10/MM2636_d N_WL<44>_XI10/MM2636_g N_BL<3>_XI10/MM2636_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2615 N_VSS_XI10/MM2615_d N_WL<43>_XI10/MM2615_g XI10/NET4860
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2792 N_VSS_XI10/MM2792_d N_WL<42>_XI10/MM2792_g N_BL<3>_XI10/MM2792_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2614 N_VSS_XI10/MM2614_d N_WL<41>_XI10/MM2614_g XI10/NET4864
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2611 N_VSS_XI10/MM2611_d N_WL<40>_XI10/MM2611_g N_BL<3>_XI10/MM2611_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2971 N_VSS_XI10/MM2971_d N_WL<39>_XI10/MM2971_g XI10/NET5380
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2928 N_VSS_XI10/MM2928_d N_WL<38>_XI10/MM2928_g N_BL<3>_XI10/MM2928_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2996 N_VSS_XI10/MM2996_d N_WL<37>_XI10/MM2996_g XI10/NET5316
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3055 N_VSS_XI10/MM3055_d N_WL<36>_XI10/MM3055_g N_BL<3>_XI10/MM3055_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3076 N_VSS_XI10/MM3076_d N_WL<35>_XI10/MM3076_g XI10/NET5112
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2899 N_VSS_XI10/MM2899_d N_WL<34>_XI10/MM2899_g N_BL<3>_XI10/MM2899_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2948 N_VSS_XI10/MM2948_d N_WL<33>_XI10/MM2948_g XI10/NET5392
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3080 N_VSS_XI10/MM3080_d N_WL<32>_XI10/MM3080_g N_BL<3>_XI10/MM3080_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1684 N_VSS_XI10/MM1684_d N_WL<31>_XI10/MM1684_g XI10/NET2200
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1739 N_VSS_XI10/MM1739_d N_WL<30>_XI10/MM1739_g N_BL<3>_XI10/MM1739_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1655 N_VSS_XI10/MM1655_d N_WL<29>_XI10/MM1655_g XI10/NET2280
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1612 N_VSS_XI10/MM1612_d N_WL<28>_XI10/MM1612_g N_BL<3>_XI10/MM1612_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1813 N_VSS_XI10/MM1813_d N_WL<27>_XI10/MM1813_g XI10/NET3004
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1768 N_VSS_XI10/MM1768_d N_WL<26>_XI10/MM1768_g N_BL<3>_XI10/MM1768_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1590 N_VSS_XI10/MM1590_d N_WL<25>_XI10/MM1590_g XI10/NET2428
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1587 N_VSS_XI10/MM1587_d N_WL<24>_XI10/MM1587_g N_BL<3>_XI10/MM1587_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1947 N_VSS_XI10/MM1947_d N_WL<23>_XI10/MM1947_g XI10/NET2768
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1904 N_VSS_XI10/MM1904_d N_WL<22>_XI10/MM1904_g N_BL<3>_XI10/MM1904_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1972 N_VSS_XI10/MM1972_d N_WL<21>_XI10/MM1972_g XI10/NET2704
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2031 N_VSS_XI10/MM2031_d N_WL<20>_XI10/MM2031_g N_BL<3>_XI10/MM2031_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1826 N_VSS_XI10/MM1826_d N_WL<19>_XI10/MM1826_g XI10/NET2960
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1875 N_VSS_XI10/MM1875_d N_WL<18>_XI10/MM1875_g N_BL<3>_XI10/MM1875_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1924 N_VSS_XI10/MM1924_d N_WL<17>_XI10/MM1924_g XI10/NET2780
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2056 N_VSS_XI10/MM2056_d N_WL<16>_XI10/MM2056_g N_BL<3>_XI10/MM2056_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1447 N_VSS_XI10/MM1447_d N_WL<15>_XI10/MM1447_g XI10/NET5696
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1392 N_VSS_XI10/MM1392_d N_WL<14>_XI10/MM1392_g N_BL<3>_XI10/MM1392_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1476 N_VSS_XI10/MM1476_d N_WL<13>_XI10/MM1476_g XI10/NET5780
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1519 N_VSS_XI10/MM1519_d N_WL<12>_XI10/MM1519_g N_BL<3>_XI10/MM1519_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1321 N_VSS_XI10/MM1321_d N_WL<11>_XI10/MM1321_g XI10/NET3432
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1363 N_VSS_XI10/MM1363_d N_WL<10>_XI10/MM1363_g N_BL<3>_XI10/MM1363_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1378 N_VSS_XI10/MM1378_d N_WL<9>_XI10/MM1378_g XI10/NET5564
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1544 N_VSS_XI10/MM1544_d N_WL<8>_XI10/MM1544_g N_BL<3>_XI10/MM1544_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1239 N_VSS_XI10/MM1239_d N_WL<7>_XI10/MM1239_g XI10/NET3152
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1185 N_VSS_XI10/MM1185_d N_WL<6>_XI10/MM1185_g N_BL<3>_XI10/MM1185_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1264 N_VSS_XI10/MM1264_d N_WL<5>_XI10/MM1264_g XI10/NET3232
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1306 N_VSS_XI10/MM1306_d N_WL<4>_XI10/MM1306_g N_BL<3>_XI10/MM1306_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1123 N_VSS_XI10/MM1123_d N_WL<3>_XI10/MM1123_g XI10/NET3416
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1178 N_VSS_XI10/MM1178_d N_WL<2>_XI10/MM1178_g N_BL<3>_XI10/MM1178_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1117 N_VSS_XI10/MM1117_d N_WL<1>_XI10/MM1117_g XI10/NET3420
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1057 N_VSS_XI10/MM1057_d N_WL<0>_XI10/MM1057_g N_BL<3>_XI10/MM1057_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2464 N_VSS_XI10/MM2464_d N_WL<63>_XI10/MM2464_g N_BL<4>_XI10/MM2464_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2422 N_VSS_XI10/MM2422_d N_WL<62>_XI10/MM2422_g XI10/NET3752
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2494 N_VSS_XI10/MM2494_d N_WL<61>_XI10/MM2494_g N_BL<4>_XI10/MM2494_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2536 N_VSS_XI10/MM2536_d N_WL<60>_XI10/MM2536_g XI10/NET5044
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2340 N_VSS_XI10/MM2340_d N_WL<59>_XI10/MM2340_g N_BL<4>_XI10/MM2340_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2380 N_VSS_XI10/MM2380_d N_WL<58>_XI10/MM2380_g XI10/NET3844
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2559 N_VSS_XI10/MM2559_d N_WL<57>_XI10/MM2559_g N_BL<4>_XI10/MM2559_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2551 N_VSS_XI10/MM2551_d N_WL<56>_XI10/MM2551_g XI10/NET4988
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2203 N_VSS_XI10/MM2203_d N_WL<55>_XI10/MM2203_g N_BL<4>_XI10/MM2203_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2244 N_VSS_XI10/MM2244_d N_WL<54>_XI10/MM2244_g XI10/NET4088
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2173 N_VSS_XI10/MM2173_d N_WL<53>_XI10/MM2173_g N_BL<4>_XI10/MM2173_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2126 N_VSS_XI10/MM2126_d N_WL<52>_XI10/MM2126_g XI10/NET3480
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2327 N_VSS_XI10/MM2327_d N_WL<51>_XI10/MM2327_g N_BL<4>_XI10/MM2327_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2282 N_VSS_XI10/MM2282_d N_WL<50>_XI10/MM2282_g XI10/NET4012
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2108 N_VSS_XI10/MM2108_d N_WL<49>_XI10/MM2108_g N_BL<4>_XI10/MM2108_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2255 N_VSS_XI10/MM2255_d N_WL<48>_XI10/MM2255_g XI10/NET4044
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2715 N_VSS_XI10/MM2715_d N_WL<47>_XI10/MM2715_g N_BL<4>_XI10/MM2715_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2756 N_VSS_XI10/MM2756_d N_WL<46>_XI10/MM2756_g XI10/NET4556
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2685 N_VSS_XI10/MM2685_d N_WL<45>_XI10/MM2685_g N_BL<4>_XI10/MM2685_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2638 N_VSS_XI10/MM2638_d N_WL<44>_XI10/MM2638_g XI10/NET4772
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2839 N_VSS_XI10/MM2839_d N_WL<43>_XI10/MM2839_g N_BL<4>_XI10/MM2839_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2794 N_VSS_XI10/MM2794_d N_WL<42>_XI10/MM2794_g XI10/NET4480
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2620 N_VSS_XI10/MM2620_d N_WL<41>_XI10/MM2620_g N_BL<4>_XI10/MM2620_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2627 N_VSS_XI10/MM2627_d N_WL<40>_XI10/MM2627_g XI10/NET4812
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2976 N_VSS_XI10/MM2976_d N_WL<39>_XI10/MM2976_g N_BL<4>_XI10/MM2976_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2930 N_VSS_XI10/MM2930_d N_WL<38>_XI10/MM2930_g XI10/NET5436
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3006 N_VSS_XI10/MM3006_d N_WL<37>_XI10/MM3006_g N_BL<4>_XI10/MM3006_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3048 N_VSS_XI10/MM3048_d N_WL<36>_XI10/MM3048_g XI10/NET5220
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2852 N_VSS_XI10/MM2852_d N_WL<35>_XI10/MM2852_g N_BL<4>_XI10/MM2852_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2892 N_VSS_XI10/MM2892_d N_WL<34>_XI10/MM2892_g XI10/NET4312
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3071 N_VSS_XI10/MM3071_d N_WL<33>_XI10/MM3071_g N_BL<4>_XI10/MM3071_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2924 N_VSS_XI10/MM2924_d N_WL<32>_XI10/MM2924_g XI10/NET5460
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1691 N_VSS_XI10/MM1691_d N_WL<31>_XI10/MM1691_g N_BL<4>_XI10/MM1691_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1732 N_VSS_XI10/MM1732_d N_WL<30>_XI10/MM1732_g XI10/NET2120
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1661 N_VSS_XI10/MM1661_d N_WL<29>_XI10/MM1661_g N_BL<4>_XI10/MM1661_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1614 N_VSS_XI10/MM1614_d N_WL<28>_XI10/MM1614_g XI10/NET2336
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1815 N_VSS_XI10/MM1815_d N_WL<27>_XI10/MM1815_g N_BL<4>_XI10/MM1815_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1770 N_VSS_XI10/MM1770_d N_WL<26>_XI10/MM1770_g XI10/NET2044
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1596 N_VSS_XI10/MM1596_d N_WL<25>_XI10/MM1596_g N_BL<4>_XI10/MM1596_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1603 N_VSS_XI10/MM1603_d N_WL<24>_XI10/MM1603_g XI10/NET2376
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1952 N_VSS_XI10/MM1952_d N_WL<23>_XI10/MM1952_g N_BL<4>_XI10/MM1952_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1906 N_VSS_XI10/MM1906_d N_WL<22>_XI10/MM1906_g XI10/NET2824
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1982 N_VSS_XI10/MM1982_d N_WL<21>_XI10/MM1982_g N_BL<4>_XI10/MM1982_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2024 N_VSS_XI10/MM2024_d N_WL<20>_XI10/MM2024_g XI10/NET02632
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1828 N_VSS_XI10/MM1828_d N_WL<19>_XI10/MM1828_g N_BL<4>_XI10/MM1828_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1868 N_VSS_XI10/MM1868_d N_WL<18>_XI10/MM1868_g XI10/NET2900
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2047 N_VSS_XI10/MM2047_d N_WL<17>_XI10/MM2047_g N_BL<4>_XI10/MM2047_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1984 N_VSS_XI10/MM1984_d N_WL<16>_XI10/MM1984_g XI10/NET2660
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1440 N_VSS_XI10/MM1440_d N_WL<15>_XI10/MM1440_g N_BL<4>_XI10/MM1440_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1399 N_VSS_XI10/MM1399_d N_WL<14>_XI10/MM1399_g XI10/NET5616
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1470 N_VSS_XI10/MM1470_d N_WL<13>_XI10/MM1470_g N_BL<4>_XI10/MM1470_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1512 N_VSS_XI10/MM1512_d N_WL<12>_XI10/MM1512_g XI10/NET1856
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1316 N_VSS_XI10/MM1316_d N_WL<11>_XI10/MM1316_g N_BL<4>_XI10/MM1316_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1361 N_VSS_XI10/MM1361_d N_WL<10>_XI10/MM1361_g XI10/NET5540
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1535 N_VSS_XI10/MM1535_d N_WL<9>_XI10/MM1535_g N_BL<4>_XI10/MM1535_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1388 N_VSS_XI10/MM1388_d N_WL<8>_XI10/MM1388_g XI10/NET5572
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1232 N_VSS_XI10/MM1232_d N_WL<7>_XI10/MM1232_g N_BL<4>_XI10/MM1232_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1192 N_VSS_XI10/MM1192_d N_WL<6>_XI10/MM1192_g XI10/NET3072
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1259 N_VSS_XI10/MM1259_d N_WL<5>_XI10/MM1259_g N_BL<4>_XI10/MM1259_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1304 N_VSS_XI10/MM1304_d N_WL<4>_XI10/MM1304_g XI10/NET3288
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1131 N_VSS_XI10/MM1131_d N_WL<3>_XI10/MM1131_g N_BL<4>_XI10/MM1131_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1176 N_VSS_XI10/MM1176_d N_WL<2>_XI10/MM1176_g XI10/NET1972
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1112 N_VSS_XI10/MM1112_d N_WL<1>_XI10/MM1112_g N_BL<4>_XI10/MM1112_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1059 N_VSS_XI10/MM1059_d N_WL<0>_XI10/MM1059_g XI10/NET3360
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI16/XI16/XI1/MM10 N_XI16/XI16/NET40_XI16/XI16/XI1/MM10_d
+ N_YOUT<5>_XI16/XI16/XI1/MM10_g N_VSS_XI16/XI16/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI15/XI1/MM10 N_XI16/XI15/NET40_XI16/XI15/XI1/MM10_d
+ N_YOUT<4>_XI16/XI15/XI1/MM10_g N_VSS_XI16/XI15/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI16/MM1 N_BL<5>_XI16/XI16/MM1_d N_XI16/XI16/NET40_XI16/XI16/MM1_g
+ N_DL<0>_XI16/XI16/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI15/MM1 N_BL<4>_XI16/XI15/MM1_d N_XI16/XI15/NET40_XI16/XI15/MM1_g
+ N_DL<0>_XI16/XI15/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2462 N_VSS_XI10/MM2462_d N_WL<63>_XI10/MM2462_g XI10/NET3700
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2417 N_VSS_XI10/MM2417_d N_WL<62>_XI10/MM2417_g N_BL<5>_XI10/MM2417_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2513 N_VSS_XI10/MM2513_d N_WL<61>_XI10/MM2513_g XI10/NET5068
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2542 N_VSS_XI10/MM2542_d N_WL<60>_XI10/MM2542_g N_BL<5>_XI10/MM2542_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2337 N_VSS_XI10/MM2337_d N_WL<59>_XI10/MM2337_g XI10/NET3908
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2386 N_VSS_XI10/MM2386_d N_WL<58>_XI10/MM2386_g N_BL<5>_XI10/MM2386_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2560 N_VSS_XI10/MM2560_d N_WL<57>_XI10/MM2560_g XI10/NET4952
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2553 N_VSS_XI10/MM2553_d N_WL<56>_XI10/MM2553_g N_BL<5>_XI10/MM2553_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2200 N_VSS_XI10/MM2200_d N_WL<55>_XI10/MM2200_g XI10/NET4156
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2250 N_VSS_XI10/MM2250_d N_WL<54>_XI10/MM2250_g N_BL<5>_XI10/MM2250_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2170 N_VSS_XI10/MM2170_d N_WL<53>_XI10/MM2170_g XI10/NET4236
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2125 N_VSS_XI10/MM2125_d N_WL<52>_XI10/MM2125_g N_BL<5>_XI10/MM2125_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2325 N_VSS_XI10/MM2325_d N_WL<51>_XI10/MM2325_g XI10/NET3948
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2281 N_VSS_XI10/MM2281_d N_WL<50>_XI10/MM2281_g N_BL<5>_XI10/MM2281_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2081 N_VSS_XI10/MM2081_d N_WL<49>_XI10/MM2081_g XI10/NET3596
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2114 N_VSS_XI10/MM2114_d N_WL<48>_XI10/MM2114_g N_BL<5>_XI10/MM2114_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2712 N_VSS_XI10/MM2712_d N_WL<47>_XI10/MM2712_g XI10/NET4624
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2762 N_VSS_XI10/MM2762_d N_WL<46>_XI10/MM2762_g N_BL<5>_XI10/MM2762_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2682 N_VSS_XI10/MM2682_d N_WL<45>_XI10/MM2682_g XI10/NET4704
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2637 N_VSS_XI10/MM2637_d N_WL<44>_XI10/MM2637_g N_BL<5>_XI10/MM2637_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2822 N_VSS_XI10/MM2822_d N_WL<43>_XI10/MM2822_g XI10/NET4436
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2793 N_VSS_XI10/MM2793_d N_WL<42>_XI10/MM2793_g N_BL<5>_XI10/MM2793_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2618 N_VSS_XI10/MM2618_d N_WL<41>_XI10/MM2618_g XI10/NET4848
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2626 N_VSS_XI10/MM2626_d N_WL<40>_XI10/MM2626_g N_BL<5>_XI10/MM2626_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2974 N_VSS_XI10/MM2974_d N_WL<39>_XI10/MM2974_g XI10/NET5368
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2929 N_VSS_XI10/MM2929_d N_WL<38>_XI10/MM2929_g N_BL<5>_XI10/MM2929_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3001 N_VSS_XI10/MM3001_d N_WL<37>_XI10/MM3001_g XI10/NET5300
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3054 N_VSS_XI10/MM3054_d N_WL<36>_XI10/MM3054_g N_BL<5>_XI10/MM3054_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2849 N_VSS_XI10/MM2849_d N_WL<35>_XI10/MM2849_g XI10/NET4376
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2898 N_VSS_XI10/MM2898_d N_WL<34>_XI10/MM2898_g N_BL<5>_XI10/MM2898_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3068 N_VSS_XI10/MM3068_d N_WL<33>_XI10/MM3068_g XI10/NET5144
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3065 N_VSS_XI10/MM3065_d N_WL<32>_XI10/MM3065_g N_BL<5>_XI10/MM3065_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1688 N_VSS_XI10/MM1688_d N_WL<31>_XI10/MM1688_g XI10/NET2188
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1738 N_VSS_XI10/MM1738_d N_WL<30>_XI10/MM1738_g N_BL<5>_XI10/MM1738_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1658 N_VSS_XI10/MM1658_d N_WL<29>_XI10/MM1658_g XI10/NET2268
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1613 N_VSS_XI10/MM1613_d N_WL<28>_XI10/MM1613_g N_BL<5>_XI10/MM1613_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1814 N_VSS_XI10/MM1814_d N_WL<27>_XI10/MM1814_g XI10/NET3000
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1769 N_VSS_XI10/MM1769_d N_WL<26>_XI10/MM1769_g N_BL<5>_XI10/MM1769_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1594 N_VSS_XI10/MM1594_d N_WL<25>_XI10/MM1594_g XI10/NET2412
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1602 N_VSS_XI10/MM1602_d N_WL<24>_XI10/MM1602_g N_BL<5>_XI10/MM1602_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1950 N_VSS_XI10/MM1950_d N_WL<23>_XI10/MM1950_g XI10/NET2756
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1905 N_VSS_XI10/MM1905_d N_WL<22>_XI10/MM1905_g N_BL<5>_XI10/MM1905_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1977 N_VSS_XI10/MM1977_d N_WL<21>_XI10/MM1977_g XI10/NET2688
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2030 N_VSS_XI10/MM2030_d N_WL<20>_XI10/MM2030_g N_BL<5>_XI10/MM2030_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1829 N_VSS_XI10/MM1829_d N_WL<19>_XI10/MM1829_g XI10/NET2948
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1874 N_VSS_XI10/MM1874_d N_WL<18>_XI10/MM1874_g N_BL<5>_XI10/MM1874_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2044 N_VSS_XI10/MM2044_d N_WL<17>_XI10/MM2044_g XI10/NET2532
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2041 N_VSS_XI10/MM2041_d N_WL<16>_XI10/MM2041_g N_BL<5>_XI10/MM2041_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1443 N_VSS_XI10/MM1443_d N_WL<15>_XI10/MM1443_g XI10/NET5684
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1393 N_VSS_XI10/MM1393_d N_WL<14>_XI10/MM1393_g N_BL<5>_XI10/MM1393_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1473 N_VSS_XI10/MM1473_d N_WL<13>_XI10/MM1473_g XI10/NET5768
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1518 N_VSS_XI10/MM1518_d N_WL<12>_XI10/MM1518_g N_BL<5>_XI10/MM1518_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1318 N_VSS_XI10/MM1318_d N_WL<11>_XI10/MM1318_g XI10/NET3356
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1362 N_VSS_XI10/MM1362_d N_WL<10>_XI10/MM1362_g N_BL<5>_XI10/MM1362_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1532 N_VSS_XI10/MM1532_d N_WL<9>_XI10/MM1532_g XI10/NET1780
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1529 N_VSS_XI10/MM1529_d N_WL<8>_XI10/MM1529_g N_BL<5>_XI10/MM1529_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1235 N_VSS_XI10/MM1235_d N_WL<7>_XI10/MM1235_g XI10/NET3140
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1186 N_VSS_XI10/MM1186_d N_WL<6>_XI10/MM1186_g N_BL<5>_XI10/MM1186_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1261 N_VSS_XI10/MM1261_d N_WL<5>_XI10/MM1261_g XI10/NET3220
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1305 N_VSS_XI10/MM1305_d N_WL<4>_XI10/MM1305_g N_BL<5>_XI10/MM1305_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1148 N_VSS_XI10/MM1148_d N_WL<3>_XI10/MM1148_g XI10/NET1928
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1177 N_VSS_XI10/MM1177_d N_WL<2>_XI10/MM1177_g N_BL<5>_XI10/MM1177_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1114 N_VSS_XI10/MM1114_d N_WL<1>_XI10/MM1114_g XI10/NET3404
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1058 N_VSS_XI10/MM1058_d N_WL<0>_XI10/MM1058_g N_BL<5>_XI10/MM1058_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2465 N_VSS_XI10/MM2465_d N_WL<63>_XI10/MM2465_g N_BL<6>_XI10/MM2465_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2415 N_VSS_XI10/MM2415_d N_WL<62>_XI10/MM2415_g XI10/NET3780
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2493 N_VSS_XI10/MM2493_d N_WL<61>_XI10/MM2493_g N_BL<6>_XI10/MM2493_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2537 N_VSS_XI10/MM2537_d N_WL<60>_XI10/MM2537_g XI10/NET5040
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2339 N_VSS_XI10/MM2339_d N_WL<59>_XI10/MM2339_g N_BL<6>_XI10/MM2339_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2381 N_VSS_XI10/MM2381_d N_WL<58>_XI10/MM2381_g XI10/NET3840
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2558 N_VSS_XI10/MM2558_d N_WL<57>_XI10/MM2558_g N_BL<6>_XI10/MM2558_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2552 N_VSS_XI10/MM2552_d N_WL<56>_XI10/MM2552_g XI10/NET4984
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2202 N_VSS_XI10/MM2202_d N_WL<55>_XI10/MM2202_g N_BL<6>_XI10/MM2202_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2245 N_VSS_XI10/MM2245_d N_WL<54>_XI10/MM2245_g XI10/NET4084
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2174 N_VSS_XI10/MM2174_d N_WL<53>_XI10/MM2174_g N_BL<6>_XI10/MM2174_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2127 N_VSS_XI10/MM2127_d N_WL<52>_XI10/MM2127_g XI10/NET3476
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2328 N_VSS_XI10/MM2328_d N_WL<51>_XI10/MM2328_g N_BL<6>_XI10/MM2328_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2283 N_VSS_XI10/MM2283_d N_WL<50>_XI10/MM2283_g XI10/NET4008
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2109 N_VSS_XI10/MM2109_d N_WL<49>_XI10/MM2109_g N_BL<6>_XI10/MM2109_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2078 N_VSS_XI10/MM2078_d N_WL<48>_XI10/MM2078_g XI10/NET3604
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2714 N_VSS_XI10/MM2714_d N_WL<47>_XI10/MM2714_g N_BL<6>_XI10/MM2714_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2757 N_VSS_XI10/MM2757_d N_WL<46>_XI10/MM2757_g XI10/NET4552
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2686 N_VSS_XI10/MM2686_d N_WL<45>_XI10/MM2686_g N_BL<6>_XI10/MM2686_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2639 N_VSS_XI10/MM2639_d N_WL<44>_XI10/MM2639_g XI10/NET4768
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2840 N_VSS_XI10/MM2840_d N_WL<43>_XI10/MM2840_g N_BL<6>_XI10/MM2840_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2795 N_VSS_XI10/MM2795_d N_WL<42>_XI10/MM2795_g XI10/NET4476
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2621 N_VSS_XI10/MM2621_d N_WL<41>_XI10/MM2621_g N_BL<6>_XI10/MM2621_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2628 N_VSS_XI10/MM2628_d N_WL<40>_XI10/MM2628_g XI10/NET4808
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2977 N_VSS_XI10/MM2977_d N_WL<39>_XI10/MM2977_g N_BL<6>_XI10/MM2977_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2931 N_VSS_XI10/MM2931_d N_WL<38>_XI10/MM2931_g XI10/NET5432
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3005 N_VSS_XI10/MM3005_d N_WL<37>_XI10/MM3005_g N_BL<6>_XI10/MM3005_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3049 N_VSS_XI10/MM3049_d N_WL<36>_XI10/MM3049_g XI10/NET5216
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2851 N_VSS_XI10/MM2851_d N_WL<35>_XI10/MM2851_g N_BL<6>_XI10/MM2851_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2893 N_VSS_XI10/MM2893_d N_WL<34>_XI10/MM2893_g XI10/NET4308
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3070 N_VSS_XI10/MM3070_d N_WL<33>_XI10/MM3070_g N_BL<6>_XI10/MM3070_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2997 N_VSS_XI10/MM2997_d N_WL<32>_XI10/MM2997_g XI10/NET5312
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1690 N_VSS_XI10/MM1690_d N_WL<31>_XI10/MM1690_g N_BL<6>_XI10/MM1690_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1733 N_VSS_XI10/MM1733_d N_WL<30>_XI10/MM1733_g XI10/NET2116
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1662 N_VSS_XI10/MM1662_d N_WL<29>_XI10/MM1662_g N_BL<6>_XI10/MM1662_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1615 N_VSS_XI10/MM1615_d N_WL<28>_XI10/MM1615_g XI10/NET2332
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1816 N_VSS_XI10/MM1816_d N_WL<27>_XI10/MM1816_g N_BL<6>_XI10/MM1816_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1771 N_VSS_XI10/MM1771_d N_WL<26>_XI10/MM1771_g XI10/NET2040
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1597 N_VSS_XI10/MM1597_d N_WL<25>_XI10/MM1597_g N_BL<6>_XI10/MM1597_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1604 N_VSS_XI10/MM1604_d N_WL<24>_XI10/MM1604_g XI10/NET2372
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1953 N_VSS_XI10/MM1953_d N_WL<23>_XI10/MM1953_g N_BL<6>_XI10/MM1953_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1907 N_VSS_XI10/MM1907_d N_WL<22>_XI10/MM1907_g XI10/NET2820
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1981 N_VSS_XI10/MM1981_d N_WL<21>_XI10/MM1981_g N_BL<6>_XI10/MM1981_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2025 N_VSS_XI10/MM2025_d N_WL<20>_XI10/MM2025_g XI10/NET02628
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1827 N_VSS_XI10/MM1827_d N_WL<19>_XI10/MM1827_g N_BL<6>_XI10/MM1827_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1869 N_VSS_XI10/MM1869_d N_WL<18>_XI10/MM1869_g XI10/NET2896
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2046 N_VSS_XI10/MM2046_d N_WL<17>_XI10/MM2046_g N_BL<6>_XI10/MM2046_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2035 N_VSS_XI10/MM2035_d N_WL<16>_XI10/MM2035_g XI10/NET2564
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1441 N_VSS_XI10/MM1441_d N_WL<15>_XI10/MM1441_g N_BL<6>_XI10/MM1441_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1398 N_VSS_XI10/MM1398_d N_WL<14>_XI10/MM1398_g XI10/NET5612
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1469 N_VSS_XI10/MM1469_d N_WL<13>_XI10/MM1469_g N_BL<6>_XI10/MM1469_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1513 N_VSS_XI10/MM1513_d N_WL<12>_XI10/MM1513_g XI10/NET1852
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1315 N_VSS_XI10/MM1315_d N_WL<11>_XI10/MM1315_g N_BL<6>_XI10/MM1315_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1360 N_VSS_XI10/MM1360_d N_WL<10>_XI10/MM1360_g XI10/NET5536
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1534 N_VSS_XI10/MM1534_d N_WL<9>_XI10/MM1534_g N_BL<6>_XI10/MM1534_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1523 N_VSS_XI10/MM1523_d N_WL<8>_XI10/MM1523_g XI10/NET1812
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1233 N_VSS_XI10/MM1233_d N_WL<7>_XI10/MM1233_g N_BL<6>_XI10/MM1233_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1191 N_VSS_XI10/MM1191_d N_WL<6>_XI10/MM1191_g XI10/NET3068
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1258 N_VSS_XI10/MM1258_d N_WL<5>_XI10/MM1258_g N_BL<6>_XI10/MM1258_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1303 N_VSS_XI10/MM1303_d N_WL<4>_XI10/MM1303_g XI10/NET3284
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1130 N_VSS_XI10/MM1130_d N_WL<3>_XI10/MM1130_g N_BL<6>_XI10/MM1130_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1175 N_VSS_XI10/MM1175_d N_WL<2>_XI10/MM1175_g XI10/NET1968
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1111 N_VSS_XI10/MM1111_d N_WL<1>_XI10/MM1111_g N_BL<6>_XI10/MM1111_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1060 N_VSS_XI10/MM1060_d N_WL<0>_XI10/MM1060_g XI10/NET3348
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI16/XI18/XI1/MM10 N_XI16/XI18/NET40_XI16/XI18/XI1/MM10_d
+ N_YOUT<7>_XI16/XI18/XI1/MM10_g N_VSS_XI16/XI18/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI17/XI1/MM10 N_XI16/XI17/NET40_XI16/XI17/XI1/MM10_d
+ N_YOUT<6>_XI16/XI17/XI1/MM10_g N_VSS_XI16/XI17/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI18/MM1 N_BL<7>_XI16/XI18/MM1_d N_XI16/XI18/NET40_XI16/XI18/MM1_g
+ N_DL<0>_XI16/XI18/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI16/XI17/MM1 N_BL<6>_XI16/XI17/MM1_d N_XI16/XI17/NET40_XI16/XI17/MM1_g
+ N_DL<0>_XI16/XI17/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2463 N_VSS_XI10/MM2463_d N_WL<63>_XI10/MM2463_g XI10/NET3696
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2420 N_VSS_XI10/MM2420_d N_WL<62>_XI10/MM2420_g N_BL<7>_XI10/MM2420_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2483 N_VSS_XI10/MM2483_d N_WL<61>_XI10/MM2483_g XI10/NET3652
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2539 N_VSS_XI10/MM2539_d N_WL<60>_XI10/MM2539_g N_BL<7>_XI10/MM2539_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2338 N_VSS_XI10/MM2338_d N_WL<59>_XI10/MM2338_g XI10/NET3904
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2383 N_VSS_XI10/MM2383_d N_WL<58>_XI10/MM2383_g N_BL<7>_XI10/MM2383_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2561 N_VSS_XI10/MM2561_d N_WL<57>_XI10/MM2561_g XI10/NET4948
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2550 N_VSS_XI10/MM2550_d N_WL<56>_XI10/MM2550_g N_BL<7>_XI10/MM2550_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2201 N_VSS_XI10/MM2201_d N_WL<55>_XI10/MM2201_g XI10/NET4152
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2247 N_VSS_XI10/MM2247_d N_WL<54>_XI10/MM2247_g N_BL<7>_XI10/MM2247_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2172 N_VSS_XI10/MM2172_d N_WL<53>_XI10/MM2172_g XI10/NET4228
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2128 N_VSS_XI10/MM2128_d N_WL<52>_XI10/MM2128_g N_BL<7>_XI10/MM2128_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2326 N_VSS_XI10/MM2326_d N_WL<51>_XI10/MM2326_g XI10/NET3944
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2284 N_VSS_XI10/MM2284_d N_WL<50>_XI10/MM2284_g N_BL<7>_XI10/MM2284_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2102 N_VSS_XI10/MM2102_d N_WL<49>_XI10/MM2102_g XI10/NET3572
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2117 N_VSS_XI10/MM2117_d N_WL<48>_XI10/MM2117_g N_BL<7>_XI10/MM2117_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2713 N_VSS_XI10/MM2713_d N_WL<47>_XI10/MM2713_g XI10/NET4620
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2759 N_VSS_XI10/MM2759_d N_WL<46>_XI10/MM2759_g N_BL<7>_XI10/MM2759_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2684 N_VSS_XI10/MM2684_d N_WL<45>_XI10/MM2684_g XI10/NET4696
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2640 N_VSS_XI10/MM2640_d N_WL<44>_XI10/MM2640_g N_BL<7>_XI10/MM2640_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2834 N_VSS_XI10/MM2834_d N_WL<43>_XI10/MM2834_g XI10/NET4428
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2796 N_VSS_XI10/MM2796_d N_WL<42>_XI10/MM2796_g N_BL<7>_XI10/MM2796_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2619 N_VSS_XI10/MM2619_d N_WL<41>_XI10/MM2619_g XI10/NET4844
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2629 N_VSS_XI10/MM2629_d N_WL<40>_XI10/MM2629_g N_BL<7>_XI10/MM2629_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2975 N_VSS_XI10/MM2975_d N_WL<39>_XI10/MM2975_g XI10/NET5364
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2932 N_VSS_XI10/MM2932_d N_WL<38>_XI10/MM2932_g N_BL<7>_XI10/MM2932_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3003 N_VSS_XI10/MM3003_d N_WL<37>_XI10/MM3003_g XI10/NET5292
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3051 N_VSS_XI10/MM3051_d N_WL<36>_XI10/MM3051_g N_BL<7>_XI10/MM3051_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2850 N_VSS_XI10/MM2850_d N_WL<35>_XI10/MM2850_g XI10/NET4372
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2895 N_VSS_XI10/MM2895_d N_WL<34>_XI10/MM2895_g N_BL<7>_XI10/MM2895_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3069 N_VSS_XI10/MM3069_d N_WL<33>_XI10/MM3069_g XI10/NET5140
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3062 N_VSS_XI10/MM3062_d N_WL<32>_XI10/MM3062_g N_BL<7>_XI10/MM3062_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1689 N_VSS_XI10/MM1689_d N_WL<31>_XI10/MM1689_g XI10/NET2184
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1735 N_VSS_XI10/MM1735_d N_WL<30>_XI10/MM1735_g N_BL<7>_XI10/MM1735_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1660 N_VSS_XI10/MM1660_d N_WL<29>_XI10/MM1660_g XI10/NET2260
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1616 N_VSS_XI10/MM1616_d N_WL<28>_XI10/MM1616_g N_BL<7>_XI10/MM1616_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1817 N_VSS_XI10/MM1817_d N_WL<27>_XI10/MM1817_g XI10/NET2988
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1772 N_VSS_XI10/MM1772_d N_WL<26>_XI10/MM1772_g N_BL<7>_XI10/MM1772_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1595 N_VSS_XI10/MM1595_d N_WL<25>_XI10/MM1595_g XI10/NET2408
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1605 N_VSS_XI10/MM1605_d N_WL<24>_XI10/MM1605_g N_BL<7>_XI10/MM1605_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1951 N_VSS_XI10/MM1951_d N_WL<23>_XI10/MM1951_g XI10/NET2752
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1908 N_VSS_XI10/MM1908_d N_WL<22>_XI10/MM1908_g N_BL<7>_XI10/MM1908_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1979 N_VSS_XI10/MM1979_d N_WL<21>_XI10/MM1979_g XI10/NET2680
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2027 N_VSS_XI10/MM2027_d N_WL<20>_XI10/MM2027_g N_BL<7>_XI10/MM2027_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1830 N_VSS_XI10/MM1830_d N_WL<19>_XI10/MM1830_g XI10/NET2944
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1871 N_VSS_XI10/MM1871_d N_WL<18>_XI10/MM1871_g N_BL<7>_XI10/MM1871_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2045 N_VSS_XI10/MM2045_d N_WL<17>_XI10/MM2045_g XI10/NET2528
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2038 N_VSS_XI10/MM2038_d N_WL<16>_XI10/MM2038_g N_BL<7>_XI10/MM2038_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1442 N_VSS_XI10/MM1442_d N_WL<15>_XI10/MM1442_g XI10/NET5680
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1396 N_VSS_XI10/MM1396_d N_WL<14>_XI10/MM1396_g N_BL<7>_XI10/MM1396_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1471 N_VSS_XI10/MM1471_d N_WL<13>_XI10/MM1471_g XI10/NET5760
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1515 N_VSS_XI10/MM1515_d N_WL<12>_XI10/MM1515_g N_BL<7>_XI10/MM1515_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1317 N_VSS_XI10/MM1317_d N_WL<11>_XI10/MM1317_g XI10/NET3352
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1359 N_VSS_XI10/MM1359_d N_WL<10>_XI10/MM1359_g N_BL<7>_XI10/MM1359_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1533 N_VSS_XI10/MM1533_d N_WL<9>_XI10/MM1533_g XI10/NET1776
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1526 N_VSS_XI10/MM1526_d N_WL<8>_XI10/MM1526_g N_BL<7>_XI10/MM1526_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1234 N_VSS_XI10/MM1234_d N_WL<7>_XI10/MM1234_g XI10/NET3136
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1189 N_VSS_XI10/MM1189_d N_WL<6>_XI10/MM1189_g N_BL<7>_XI10/MM1189_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1260 N_VSS_XI10/MM1260_d N_WL<5>_XI10/MM1260_g XI10/NET3212
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1302 N_VSS_XI10/MM1302_d N_WL<4>_XI10/MM1302_g N_BL<7>_XI10/MM1302_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1136 N_VSS_XI10/MM1136_d N_WL<3>_XI10/MM1136_g XI10/NET1920
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1174 N_VSS_XI10/MM1174_d N_WL<2>_XI10/MM1174_g N_BL<7>_XI10/MM1174_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1113 N_VSS_XI10/MM1113_d N_WL<1>_XI10/MM1113_g XI10/NET3400
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1061 N_VSS_XI10/MM1061_d N_WL<0>_XI10/MM1061_g N_BL<7>_XI10/MM1061_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2468 N_VSS_XI10/MM2468_d N_WL<63>_XI10/MM2468_g N_BL<8>_XI10/MM2468_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2423 N_VSS_XI10/MM2423_d N_WL<62>_XI10/MM2423_g XI10/NET3748
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2488 N_VSS_XI10/MM2488_d N_WL<61>_XI10/MM2488_g N_BL<8>_XI10/MM2488_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2540 N_VSS_XI10/MM2540_d N_WL<60>_XI10/MM2540_g XI10/NET5028
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2336 N_VSS_XI10/MM2336_d N_WL<59>_XI10/MM2336_g N_BL<8>_XI10/MM2336_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2384 N_VSS_XI10/MM2384_d N_WL<58>_XI10/MM2384_g XI10/NET3828
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2555 N_VSS_XI10/MM2555_d N_WL<57>_XI10/MM2555_g N_BL<8>_XI10/MM2555_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2573 N_VSS_XI10/MM2573_d N_WL<56>_XI10/MM2573_g XI10/NET4916
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2199 N_VSS_XI10/MM2199_d N_WL<55>_XI10/MM2199_g N_BL<8>_XI10/MM2199_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2248 N_VSS_XI10/MM2248_d N_WL<54>_XI10/MM2248_g XI10/NET4072
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2179 N_VSS_XI10/MM2179_d N_WL<53>_XI10/MM2179_g N_BL<8>_XI10/MM2179_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2130 N_VSS_XI10/MM2130_d N_WL<52>_XI10/MM2130_g XI10/NET3464
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2331 N_VSS_XI10/MM2331_d N_WL<51>_XI10/MM2331_g N_BL<8>_XI10/MM2331_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2286 N_VSS_XI10/MM2286_d N_WL<50>_XI10/MM2286_g XI10/NET3996
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2112 N_VSS_XI10/MM2112_d N_WL<49>_XI10/MM2112_g N_BL<8>_XI10/MM2112_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2094 N_VSS_XI10/MM2094_d N_WL<48>_XI10/MM2094_g XI10/NET3588
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2711 N_VSS_XI10/MM2711_d N_WL<47>_XI10/MM2711_g N_BL<8>_XI10/MM2711_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2760 N_VSS_XI10/MM2760_d N_WL<46>_XI10/MM2760_g XI10/NET4540
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2691 N_VSS_XI10/MM2691_d N_WL<45>_XI10/MM2691_g N_BL<8>_XI10/MM2691_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2642 N_VSS_XI10/MM2642_d N_WL<44>_XI10/MM2642_g XI10/NET4756
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2843 N_VSS_XI10/MM2843_d N_WL<43>_XI10/MM2843_g N_BL<8>_XI10/MM2843_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2798 N_VSS_XI10/MM2798_d N_WL<42>_XI10/MM2798_g XI10/NET4464
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2624 N_VSS_XI10/MM2624_d N_WL<41>_XI10/MM2624_g N_BL<8>_XI10/MM2624_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2632 N_VSS_XI10/MM2632_d N_WL<40>_XI10/MM2632_g XI10/NET4796
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2980 N_VSS_XI10/MM2980_d N_WL<39>_XI10/MM2980_g N_BL<8>_XI10/MM2980_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2934 N_VSS_XI10/MM2934_d N_WL<38>_XI10/MM2934_g XI10/NET5420
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3000 N_VSS_XI10/MM3000_d N_WL<37>_XI10/MM3000_g N_BL<8>_XI10/MM3000_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3052 N_VSS_XI10/MM3052_d N_WL<36>_XI10/MM3052_g XI10/NET5204
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2848 N_VSS_XI10/MM2848_d N_WL<35>_XI10/MM2848_g N_BL<8>_XI10/MM2848_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2896 N_VSS_XI10/MM2896_d N_WL<34>_XI10/MM2896_g XI10/NET4296
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3067 N_VSS_XI10/MM3067_d N_WL<33>_XI10/MM3067_g N_BL<8>_XI10/MM3067_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3008 N_VSS_XI10/MM3008_d N_WL<32>_XI10/MM3008_g XI10/NET5272
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1687 N_VSS_XI10/MM1687_d N_WL<31>_XI10/MM1687_g N_BL<8>_XI10/MM1687_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1736 N_VSS_XI10/MM1736_d N_WL<30>_XI10/MM1736_g XI10/NET2104
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1667 N_VSS_XI10/MM1667_d N_WL<29>_XI10/MM1667_g N_BL<8>_XI10/MM1667_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1618 N_VSS_XI10/MM1618_d N_WL<28>_XI10/MM1618_g XI10/NET2320
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1819 N_VSS_XI10/MM1819_d N_WL<27>_XI10/MM1819_g N_BL<8>_XI10/MM1819_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1774 N_VSS_XI10/MM1774_d N_WL<26>_XI10/MM1774_g XI10/NET2028
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1600 N_VSS_XI10/MM1600_d N_WL<25>_XI10/MM1600_g N_BL<8>_XI10/MM1600_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1608 N_VSS_XI10/MM1608_d N_WL<24>_XI10/MM1608_g XI10/NET2360
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1956 N_VSS_XI10/MM1956_d N_WL<23>_XI10/MM1956_g N_BL<8>_XI10/MM1956_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1910 N_VSS_XI10/MM1910_d N_WL<22>_XI10/MM1910_g XI10/NET2808
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1976 N_VSS_XI10/MM1976_d N_WL<21>_XI10/MM1976_g N_BL<8>_XI10/MM1976_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2028 N_VSS_XI10/MM2028_d N_WL<20>_XI10/MM2028_g XI10/NET02616
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1824 N_VSS_XI10/MM1824_d N_WL<19>_XI10/MM1824_g N_BL<8>_XI10/MM1824_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1872 N_VSS_XI10/MM1872_d N_WL<18>_XI10/MM1872_g XI10/NET2884
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2043 N_VSS_XI10/MM2043_d N_WL<17>_XI10/MM2043_g N_BL<8>_XI10/MM2043_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2039 N_VSS_XI10/MM2039_d N_WL<16>_XI10/MM2039_g XI10/NET2552
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1444 N_VSS_XI10/MM1444_d N_WL<15>_XI10/MM1444_g N_BL<8>_XI10/MM1444_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1395 N_VSS_XI10/MM1395_d N_WL<14>_XI10/MM1395_g XI10/NET5600
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1464 N_VSS_XI10/MM1464_d N_WL<13>_XI10/MM1464_g N_BL<8>_XI10/MM1464_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1516 N_VSS_XI10/MM1516_d N_WL<12>_XI10/MM1516_g XI10/NET1840
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1312 N_VSS_XI10/MM1312_d N_WL<11>_XI10/MM1312_g N_BL<8>_XI10/MM1312_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1357 N_VSS_XI10/MM1357_d N_WL<10>_XI10/MM1357_g XI10/NET5524
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1531 N_VSS_XI10/MM1531_d N_WL<9>_XI10/MM1531_g N_BL<8>_XI10/MM1531_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1527 N_VSS_XI10/MM1527_d N_WL<8>_XI10/MM1527_g XI10/NET1800
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1236 N_VSS_XI10/MM1236_d N_WL<7>_XI10/MM1236_g N_BL<8>_XI10/MM1236_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1188 N_VSS_XI10/MM1188_d N_WL<6>_XI10/MM1188_g XI10/NET3056
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1255 N_VSS_XI10/MM1255_d N_WL<5>_XI10/MM1255_g N_BL<8>_XI10/MM1255_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1300 N_VSS_XI10/MM1300_d N_WL<4>_XI10/MM1300_g XI10/NET3272
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1127 N_VSS_XI10/MM1127_d N_WL<3>_XI10/MM1127_g N_BL<8>_XI10/MM1127_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1172 N_VSS_XI10/MM1172_d N_WL<2>_XI10/MM1172_g XI10/NET1956
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1108 N_VSS_XI10/MM1108_d N_WL<1>_XI10/MM1108_g N_BL<8>_XI10/MM1108_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1063 N_VSS_XI10/MM1063_d N_WL<0>_XI10/MM1063_g XI10/NET3336
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI17/XI21/XI1/MM10 N_XI17/XI21/NET40_XI17/XI21/XI1/MM10_d
+ N_YOUT<1>_XI17/XI21/XI1/MM10_g N_VSS_XI17/XI21/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI22/XI1/MM10 N_XI17/XI22/NET40_XI17/XI22/XI1/MM10_d
+ N_YOUT<0>_XI17/XI22/XI1/MM10_g N_VSS_XI17/XI22/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI21/MM1 N_BL<9>_XI17/XI21/MM1_d N_XI17/XI21/NET40_XI17/XI21/MM1_g
+ N_DL<1>_XI17/XI21/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI22/MM1 N_BL<8>_XI17/XI22/MM1_d N_XI17/XI22/NET40_XI17/XI22/MM1_g
+ N_DL<1>_XI17/XI22/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2466 N_VSS_XI10/MM2466_d N_WL<63>_XI10/MM2466_g XI10/NET3684
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2421 N_VSS_XI10/MM2421_d N_WL<62>_XI10/MM2421_g N_BL<9>_XI10/MM2421_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2484 N_VSS_XI10/MM2484_d N_WL<61>_XI10/MM2484_g XI10/NET3648
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2538 N_VSS_XI10/MM2538_d N_WL<60>_XI10/MM2538_g N_BL<9>_XI10/MM2538_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2341 N_VSS_XI10/MM2341_d N_WL<59>_XI10/MM2341_g XI10/NET3892
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2382 N_VSS_XI10/MM2382_d N_WL<58>_XI10/MM2382_g N_BL<9>_XI10/MM2382_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2565 N_VSS_XI10/MM2565_d N_WL<57>_XI10/MM2565_g XI10/NET4932
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2548 N_VSS_XI10/MM2548_d N_WL<56>_XI10/MM2548_g N_BL<9>_XI10/MM2548_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2204 N_VSS_XI10/MM2204_d N_WL<55>_XI10/MM2204_g XI10/NET4140
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2246 N_VSS_XI10/MM2246_d N_WL<54>_XI10/MM2246_g N_BL<9>_XI10/MM2246_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2176 N_VSS_XI10/MM2176_d N_WL<53>_XI10/MM2176_g XI10/NET4212
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2129 N_VSS_XI10/MM2129_d N_WL<52>_XI10/MM2129_g N_BL<9>_XI10/MM2129_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2329 N_VSS_XI10/MM2329_d N_WL<51>_XI10/MM2329_g XI10/NET3932
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2285 N_VSS_XI10/MM2285_d N_WL<50>_XI10/MM2285_g N_BL<9>_XI10/MM2285_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2106 N_VSS_XI10/MM2106_d N_WL<49>_XI10/MM2106_g XI10/NET3556
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2119 N_VSS_XI10/MM2119_d N_WL<48>_XI10/MM2119_g N_BL<9>_XI10/MM2119_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2716 N_VSS_XI10/MM2716_d N_WL<47>_XI10/MM2716_g XI10/NET4608
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2758 N_VSS_XI10/MM2758_d N_WL<46>_XI10/MM2758_g N_BL<9>_XI10/MM2758_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2688 N_VSS_XI10/MM2688_d N_WL<45>_XI10/MM2688_g XI10/NET4680
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2641 N_VSS_XI10/MM2641_d N_WL<44>_XI10/MM2641_g N_BL<9>_XI10/MM2641_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2837 N_VSS_XI10/MM2837_d N_WL<43>_XI10/MM2837_g XI10/NET4416
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2797 N_VSS_XI10/MM2797_d N_WL<42>_XI10/MM2797_g N_BL<9>_XI10/MM2797_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2622 N_VSS_XI10/MM2622_d N_WL<41>_XI10/MM2622_g XI10/NET4832
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2631 N_VSS_XI10/MM2631_d N_WL<40>_XI10/MM2631_g N_BL<9>_XI10/MM2631_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2978 N_VSS_XI10/MM2978_d N_WL<39>_XI10/MM2978_g XI10/NET5352
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2933 N_VSS_XI10/MM2933_d N_WL<38>_XI10/MM2933_g N_BL<9>_XI10/MM2933_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3007 N_VSS_XI10/MM3007_d N_WL<37>_XI10/MM3007_g XI10/NET5276
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3050 N_VSS_XI10/MM3050_d N_WL<36>_XI10/MM3050_g N_BL<9>_XI10/MM3050_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2853 N_VSS_XI10/MM2853_d N_WL<35>_XI10/MM2853_g XI10/NET4360
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2894 N_VSS_XI10/MM2894_d N_WL<34>_XI10/MM2894_g N_BL<9>_XI10/MM2894_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3072 N_VSS_XI10/MM3072_d N_WL<33>_XI10/MM3072_g XI10/NET5128
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3060 N_VSS_XI10/MM3060_d N_WL<32>_XI10/MM3060_g N_BL<9>_XI10/MM3060_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1692 N_VSS_XI10/MM1692_d N_WL<31>_XI10/MM1692_g XI10/NET2172
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1734 N_VSS_XI10/MM1734_d N_WL<30>_XI10/MM1734_g N_BL<9>_XI10/MM1734_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1664 N_VSS_XI10/MM1664_d N_WL<29>_XI10/MM1664_g XI10/NET2244
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1617 N_VSS_XI10/MM1617_d N_WL<28>_XI10/MM1617_g N_BL<9>_XI10/MM1617_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1818 N_VSS_XI10/MM1818_d N_WL<27>_XI10/MM1818_g XI10/NET2984
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1773 N_VSS_XI10/MM1773_d N_WL<26>_XI10/MM1773_g N_BL<9>_XI10/MM1773_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1598 N_VSS_XI10/MM1598_d N_WL<25>_XI10/MM1598_g XI10/NET2396
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1607 N_VSS_XI10/MM1607_d N_WL<24>_XI10/MM1607_g N_BL<9>_XI10/MM1607_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1954 N_VSS_XI10/MM1954_d N_WL<23>_XI10/MM1954_g XI10/NET2740
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1909 N_VSS_XI10/MM1909_d N_WL<22>_XI10/MM1909_g N_BL<9>_XI10/MM1909_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1983 N_VSS_XI10/MM1983_d N_WL<21>_XI10/MM1983_g XI10/NET2664
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2026 N_VSS_XI10/MM2026_d N_WL<20>_XI10/MM2026_g N_BL<9>_XI10/MM2026_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1833 N_VSS_XI10/MM1833_d N_WL<19>_XI10/MM1833_g XI10/NET2932
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1870 N_VSS_XI10/MM1870_d N_WL<18>_XI10/MM1870_g N_BL<9>_XI10/MM1870_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2048 N_VSS_XI10/MM2048_d N_WL<17>_XI10/MM2048_g XI10/NET2516
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2036 N_VSS_XI10/MM2036_d N_WL<16>_XI10/MM2036_g N_BL<9>_XI10/MM2036_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1439 N_VSS_XI10/MM1439_d N_WL<15>_XI10/MM1439_g XI10/NET5668
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1397 N_VSS_XI10/MM1397_d N_WL<14>_XI10/MM1397_g N_BL<9>_XI10/MM1397_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1467 N_VSS_XI10/MM1467_d N_WL<13>_XI10/MM1467_g XI10/NET5744
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1514 N_VSS_XI10/MM1514_d N_WL<12>_XI10/MM1514_g N_BL<9>_XI10/MM1514_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1314 N_VSS_XI10/MM1314_d N_WL<11>_XI10/MM1314_g XI10/NET3324
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1358 N_VSS_XI10/MM1358_d N_WL<10>_XI10/MM1358_g N_BL<9>_XI10/MM1358_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1536 N_VSS_XI10/MM1536_d N_WL<9>_XI10/MM1536_g XI10/NET1764
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1524 N_VSS_XI10/MM1524_d N_WL<8>_XI10/MM1524_g N_BL<9>_XI10/MM1524_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1231 N_VSS_XI10/MM1231_d N_WL<7>_XI10/MM1231_g XI10/NET3124
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1190 N_VSS_XI10/MM1190_d N_WL<6>_XI10/MM1190_g N_BL<9>_XI10/MM1190_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1257 N_VSS_XI10/MM1257_d N_WL<5>_XI10/MM1257_g XI10/NET3196
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1301 N_VSS_XI10/MM1301_d N_WL<4>_XI10/MM1301_g N_BL<9>_XI10/MM1301_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1133 N_VSS_XI10/MM1133_d N_WL<3>_XI10/MM1133_g XI10/NET1908
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1173 N_VSS_XI10/MM1173_d N_WL<2>_XI10/MM1173_g N_BL<9>_XI10/MM1173_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1110 N_VSS_XI10/MM1110_d N_WL<1>_XI10/MM1110_g XI10/NET3388
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1062 N_VSS_XI10/MM1062_d N_WL<0>_XI10/MM1062_g N_BL<9>_XI10/MM1062_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2469 N_VSS_XI10/MM2469_d N_WL<63>_XI10/MM2469_g N_BL<10>_XI10/MM2469_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2419 N_VSS_XI10/MM2419_d N_WL<62>_XI10/MM2419_g XI10/NET3764
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2487 N_VSS_XI10/MM2487_d N_WL<61>_XI10/MM2487_g N_BL<10>_XI10/MM2487_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2541 N_VSS_XI10/MM2541_d N_WL<60>_XI10/MM2541_g XI10/NET5024
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2566 N_VSS_XI10/MM2566_d N_WL<59>_XI10/MM2566_g N_BL<10>_XI10/MM2566_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2385 N_VSS_XI10/MM2385_d N_WL<58>_XI10/MM2385_g XI10/NET3824
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2554 N_VSS_XI10/MM2554_d N_WL<57>_XI10/MM2554_g N_BL<10>_XI10/MM2554_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2589 N_VSS_XI10/MM2589_d N_WL<56>_XI10/MM2589_g XI10/NET4900
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2198 N_VSS_XI10/MM2198_d N_WL<55>_XI10/MM2198_g N_BL<10>_XI10/MM2198_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2249 N_VSS_XI10/MM2249_d N_WL<54>_XI10/MM2249_g XI10/NET4068
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2180 N_VSS_XI10/MM2180_d N_WL<53>_XI10/MM2180_g N_BL<10>_XI10/MM2180_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2131 N_VSS_XI10/MM2131_d N_WL<52>_XI10/MM2131_g XI10/NET3460
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2101 N_VSS_XI10/MM2101_d N_WL<51>_XI10/MM2101_g N_BL<10>_XI10/MM2101_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2287 N_VSS_XI10/MM2287_d N_WL<50>_XI10/MM2287_g XI10/NET3992
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2113 N_VSS_XI10/MM2113_d N_WL<49>_XI10/MM2113_g N_BL<10>_XI10/MM2113_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2115 N_VSS_XI10/MM2115_d N_WL<48>_XI10/MM2115_g XI10/NET3520
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2710 N_VSS_XI10/MM2710_d N_WL<47>_XI10/MM2710_g N_BL<10>_XI10/MM2710_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2761 N_VSS_XI10/MM2761_d N_WL<46>_XI10/MM2761_g XI10/NET4536
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2692 N_VSS_XI10/MM2692_d N_WL<45>_XI10/MM2692_g N_BL<10>_XI10/MM2692_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2643 N_VSS_XI10/MM2643_d N_WL<44>_XI10/MM2643_g XI10/NET4752
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2613 N_VSS_XI10/MM2613_d N_WL<43>_XI10/MM2613_g N_BL<10>_XI10/MM2613_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2799 N_VSS_XI10/MM2799_d N_WL<42>_XI10/MM2799_g XI10/NET4460
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2625 N_VSS_XI10/MM2625_d N_WL<41>_XI10/MM2625_g N_BL<10>_XI10/MM2625_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2683 N_VSS_XI10/MM2683_d N_WL<40>_XI10/MM2683_g XI10/NET4700
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2981 N_VSS_XI10/MM2981_d N_WL<39>_XI10/MM2981_g N_BL<10>_XI10/MM2981_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2935 N_VSS_XI10/MM2935_d N_WL<38>_XI10/MM2935_g XI10/NET5416
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2999 N_VSS_XI10/MM2999_d N_WL<37>_XI10/MM2999_g N_BL<10>_XI10/MM2999_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3053 N_VSS_XI10/MM3053_d N_WL<36>_XI10/MM3053_g XI10/NET5200
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3078 N_VSS_XI10/MM3078_d N_WL<35>_XI10/MM3078_g N_BL<10>_XI10/MM3078_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2897 N_VSS_XI10/MM2897_d N_WL<34>_XI10/MM2897_g XI10/NET4292
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3066 N_VSS_XI10/MM3066_d N_WL<33>_XI10/MM3066_g N_BL<10>_XI10/MM3066_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3059 N_VSS_XI10/MM3059_d N_WL<32>_XI10/MM3059_g XI10/NET5176
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1686 N_VSS_XI10/MM1686_d N_WL<31>_XI10/MM1686_g N_BL<10>_XI10/MM1686_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1737 N_VSS_XI10/MM1737_d N_WL<30>_XI10/MM1737_g XI10/NET2100
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1668 N_VSS_XI10/MM1668_d N_WL<29>_XI10/MM1668_g N_BL<10>_XI10/MM1668_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1619 N_VSS_XI10/MM1619_d N_WL<28>_XI10/MM1619_g XI10/NET2316
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1589 N_VSS_XI10/MM1589_d N_WL<27>_XI10/MM1589_g N_BL<10>_XI10/MM1589_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1775 N_VSS_XI10/MM1775_d N_WL<26>_XI10/MM1775_g XI10/NET2024
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1601 N_VSS_XI10/MM1601_d N_WL<25>_XI10/MM1601_g N_BL<10>_XI10/MM1601_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1659 N_VSS_XI10/MM1659_d N_WL<24>_XI10/MM1659_g XI10/NET2264
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1957 N_VSS_XI10/MM1957_d N_WL<23>_XI10/MM1957_g N_BL<10>_XI10/MM1957_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1911 N_VSS_XI10/MM1911_d N_WL<22>_XI10/MM1911_g XI10/NET2804
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1975 N_VSS_XI10/MM1975_d N_WL<21>_XI10/MM1975_g N_BL<10>_XI10/MM1975_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2029 N_VSS_XI10/MM2029_d N_WL<20>_XI10/MM2029_g XI10/NET02612
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2054 N_VSS_XI10/MM2054_d N_WL<19>_XI10/MM2054_g N_BL<10>_XI10/MM2054_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1873 N_VSS_XI10/MM1873_d N_WL<18>_XI10/MM1873_g XI10/NET2880
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2042 N_VSS_XI10/MM2042_d N_WL<17>_XI10/MM2042_g N_BL<10>_XI10/MM2042_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2040 N_VSS_XI10/MM2040_d N_WL<16>_XI10/MM2040_g XI10/NET2548
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1445 N_VSS_XI10/MM1445_d N_WL<15>_XI10/MM1445_g N_BL<10>_XI10/MM1445_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1394 N_VSS_XI10/MM1394_d N_WL<14>_XI10/MM1394_g XI10/NET5596
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1463 N_VSS_XI10/MM1463_d N_WL<13>_XI10/MM1463_g N_BL<10>_XI10/MM1463_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1517 N_VSS_XI10/MM1517_d N_WL<12>_XI10/MM1517_g XI10/NET1836
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1542 N_VSS_XI10/MM1542_d N_WL<11>_XI10/MM1542_g N_BL<10>_XI10/MM1542_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1356 N_VSS_XI10/MM1356_d N_WL<10>_XI10/MM1356_g XI10/NET5520
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1530 N_VSS_XI10/MM1530_d N_WL<9>_XI10/MM1530_g N_BL<10>_XI10/MM1530_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1528 N_VSS_XI10/MM1528_d N_WL<8>_XI10/MM1528_g XI10/NET1796
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1237 N_VSS_XI10/MM1237_d N_WL<7>_XI10/MM1237_g N_BL<10>_XI10/MM1237_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1187 N_VSS_XI10/MM1187_d N_WL<6>_XI10/MM1187_g XI10/NET3052
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1254 N_VSS_XI10/MM1254_d N_WL<5>_XI10/MM1254_g N_BL<10>_XI10/MM1254_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1299 N_VSS_XI10/MM1299_d N_WL<4>_XI10/MM1299_g XI10/NET3268
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1126 N_VSS_XI10/MM1126_d N_WL<3>_XI10/MM1126_g N_BL<10>_XI10/MM1126_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1171 N_VSS_XI10/MM1171_d N_WL<2>_XI10/MM1171_g XI10/NET1952
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1107 N_VSS_XI10/MM1107_d N_WL<1>_XI10/MM1107_g N_BL<10>_XI10/MM1107_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1064 N_VSS_XI10/MM1064_d N_WL<0>_XI10/MM1064_g XI10/NET3216
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI17/XI19/XI1/MM10 N_XI17/XI19/NET40_XI17/XI19/XI1/MM10_d
+ N_YOUT<3>_XI17/XI19/XI1/MM10_g N_VSS_XI17/XI19/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI20/XI1/MM10 N_XI17/XI20/NET40_XI17/XI20/XI1/MM10_d
+ N_YOUT<2>_XI17/XI20/XI1/MM10_g N_VSS_XI17/XI20/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI19/MM1 N_BL<11>_XI17/XI19/MM1_d N_XI17/XI19/NET40_XI17/XI19/MM1_g
+ N_DL<1>_XI17/XI19/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI20/MM1 N_BL<10>_XI17/XI20/MM1_d N_XI17/XI20/NET40_XI17/XI20/MM1_g
+ N_DL<1>_XI17/XI20/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2467 N_VSS_XI10/MM2467_d N_WL<63>_XI10/MM2467_g XI10/NET3680
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2424 N_VSS_XI10/MM2424_d N_WL<62>_XI10/MM2424_g N_BL<11>_XI10/MM2424_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2489 N_VSS_XI10/MM2489_d N_WL<61>_XI10/MM2489_g XI10/NET3632
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2535 N_VSS_XI10/MM2535_d N_WL<60>_XI10/MM2535_g N_BL<11>_XI10/MM2535_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2342 N_VSS_XI10/MM2342_d N_WL<59>_XI10/MM2342_g XI10/NET3888
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2379 N_VSS_XI10/MM2379_d N_WL<58>_XI10/MM2379_g N_BL<11>_XI10/MM2379_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2586 N_VSS_XI10/MM2586_d N_WL<57>_XI10/MM2586_g XI10/NET4908
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2492 N_VSS_XI10/MM2492_d N_WL<56>_XI10/MM2492_g N_BL<11>_XI10/MM2492_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2205 N_VSS_XI10/MM2205_d N_WL<55>_XI10/MM2205_g XI10/NET4136
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2243 N_VSS_XI10/MM2243_d N_WL<54>_XI10/MM2243_g N_BL<11>_XI10/MM2243_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2178 N_VSS_XI10/MM2178_d N_WL<53>_XI10/MM2178_g XI10/NET4204
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2132 N_VSS_XI10/MM2132_d N_WL<52>_XI10/MM2132_g N_BL<11>_XI10/MM2132_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2330 N_VSS_XI10/MM2330_d N_WL<51>_XI10/MM2330_g XI10/NET3928
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2288 N_VSS_XI10/MM2288_d N_WL<50>_XI10/MM2288_g N_BL<11>_XI10/MM2288_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2107 N_VSS_XI10/MM2107_d N_WL<49>_XI10/MM2107_g XI10/NET3552
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2175 N_VSS_XI10/MM2175_d N_WL<48>_XI10/MM2175_g N_BL<11>_XI10/MM2175_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2717 N_VSS_XI10/MM2717_d N_WL<47>_XI10/MM2717_g XI10/NET4604
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2755 N_VSS_XI10/MM2755_d N_WL<46>_XI10/MM2755_g N_BL<11>_XI10/MM2755_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2690 N_VSS_XI10/MM2690_d N_WL<45>_XI10/MM2690_g XI10/NET4672
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2644 N_VSS_XI10/MM2644_d N_WL<44>_XI10/MM2644_g N_BL<11>_XI10/MM2644_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2838 N_VSS_XI10/MM2838_d N_WL<43>_XI10/MM2838_g XI10/NET4412
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2800 N_VSS_XI10/MM2800_d N_WL<42>_XI10/MM2800_g N_BL<11>_XI10/MM2800_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2623 N_VSS_XI10/MM2623_d N_WL<41>_XI10/MM2623_g XI10/NET4828
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2687 N_VSS_XI10/MM2687_d N_WL<40>_XI10/MM2687_g N_BL<11>_XI10/MM2687_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2979 N_VSS_XI10/MM2979_d N_WL<39>_XI10/MM2979_g XI10/NET5348
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2936 N_VSS_XI10/MM2936_d N_WL<38>_XI10/MM2936_g N_BL<11>_XI10/MM2936_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3009 N_VSS_XI10/MM3009_d N_WL<37>_XI10/MM3009_g XI10/NET5268
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3047 N_VSS_XI10/MM3047_d N_WL<36>_XI10/MM3047_g N_BL<11>_XI10/MM3047_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2854 N_VSS_XI10/MM2854_d N_WL<35>_XI10/MM2854_g XI10/NET4356
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2891 N_VSS_XI10/MM2891_d N_WL<34>_XI10/MM2891_g N_BL<11>_XI10/MM2891_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3073 N_VSS_XI10/MM3073_d N_WL<33>_XI10/MM3073_g XI10/NET5124
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3004 N_VSS_XI10/MM3004_d N_WL<32>_XI10/MM3004_g N_BL<11>_XI10/MM3004_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1693 N_VSS_XI10/MM1693_d N_WL<31>_XI10/MM1693_g XI10/NET2168
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1731 N_VSS_XI10/MM1731_d N_WL<30>_XI10/MM1731_g N_BL<11>_XI10/MM1731_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1666 N_VSS_XI10/MM1666_d N_WL<29>_XI10/MM1666_g XI10/NET2236
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1620 N_VSS_XI10/MM1620_d N_WL<28>_XI10/MM1620_g N_BL<11>_XI10/MM1620_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1585 N_VSS_XI10/MM1585_d N_WL<27>_XI10/MM1585_g XI10/NET2440
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1776 N_VSS_XI10/MM1776_d N_WL<26>_XI10/MM1776_g N_BL<11>_XI10/MM1776_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1599 N_VSS_XI10/MM1599_d N_WL<25>_XI10/MM1599_g XI10/NET2392
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1663 N_VSS_XI10/MM1663_d N_WL<24>_XI10/MM1663_g N_BL<11>_XI10/MM1663_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1955 N_VSS_XI10/MM1955_d N_WL<23>_XI10/MM1955_g XI10/NET2736
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1912 N_VSS_XI10/MM1912_d N_WL<22>_XI10/MM1912_g N_BL<11>_XI10/MM1912_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1985 N_VSS_XI10/MM1985_d N_WL<21>_XI10/MM1985_g XI10/NET2656
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2023 N_VSS_XI10/MM2023_d N_WL<20>_XI10/MM2023_g N_BL<11>_XI10/MM2023_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1845 N_VSS_XI10/MM1845_d N_WL<19>_XI10/MM1845_g XI10/NET2924
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1867 N_VSS_XI10/MM1867_d N_WL<18>_XI10/MM1867_g N_BL<11>_XI10/MM1867_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2049 N_VSS_XI10/MM2049_d N_WL<17>_XI10/MM2049_g XI10/NET2512
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1980 N_VSS_XI10/MM1980_d N_WL<16>_XI10/MM1980_g N_BL<11>_XI10/MM1980_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1438 N_VSS_XI10/MM1438_d N_WL<15>_XI10/MM1438_g XI10/NET5664
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1400 N_VSS_XI10/MM1400_d N_WL<14>_XI10/MM1400_g N_BL<11>_XI10/MM1400_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1465 N_VSS_XI10/MM1465_d N_WL<13>_XI10/MM1465_g XI10/NET5736
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1511 N_VSS_XI10/MM1511_d N_WL<12>_XI10/MM1511_g N_BL<11>_XI10/MM1511_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1313 N_VSS_XI10/MM1313_d N_WL<11>_XI10/MM1313_g XI10/NET3320
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1355 N_VSS_XI10/MM1355_d N_WL<10>_XI10/MM1355_g N_BL<11>_XI10/MM1355_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1537 N_VSS_XI10/MM1537_d N_WL<9>_XI10/MM1537_g XI10/NET1760
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1468 N_VSS_XI10/MM1468_d N_WL<8>_XI10/MM1468_g N_BL<11>_XI10/MM1468_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1230 N_VSS_XI10/MM1230_d N_WL<7>_XI10/MM1230_g XI10/NET3120
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1193 N_VSS_XI10/MM1193_d N_WL<6>_XI10/MM1193_g N_BL<11>_XI10/MM1193_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1256 N_VSS_XI10/MM1256_d N_WL<5>_XI10/MM1256_g XI10/NET3188
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1298 N_VSS_XI10/MM1298_d N_WL<4>_XI10/MM1298_g N_BL<11>_XI10/MM1298_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1132 N_VSS_XI10/MM1132_d N_WL<3>_XI10/MM1132_g XI10/NET1904
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1170 N_VSS_XI10/MM1170_d N_WL<2>_XI10/MM1170_g N_BL<11>_XI10/MM1170_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1109 N_VSS_XI10/MM1109_d N_WL<1>_XI10/MM1109_g XI10/NET3384
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1065 N_VSS_XI10/MM1065_d N_WL<0>_XI10/MM1065_g N_BL<11>_XI10/MM1065_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2451 N_VSS_XI10/MM2451_d N_WL<63>_XI10/MM2451_g N_BL<12>_XI10/MM2451_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2426 N_VSS_XI10/MM2426_d N_WL<62>_XI10/MM2426_g XI10/NET3736
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2509 N_VSS_XI10/MM2509_d N_WL<61>_XI10/MM2509_g N_BL<12>_XI10/MM2509_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2544 N_VSS_XI10/MM2544_d N_WL<60>_XI10/MM2544_g XI10/NET5012
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2353 N_VSS_XI10/MM2353_d N_WL<59>_XI10/MM2353_g N_BL<12>_XI10/MM2353_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2388 N_VSS_XI10/MM2388_d N_WL<58>_XI10/MM2388_g XI10/NET3812
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2582 N_VSS_XI10/MM2582_d N_WL<57>_XI10/MM2582_g N_BL<12>_XI10/MM2582_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2412 N_VSS_XI10/MM2412_d N_WL<56>_XI10/MM2412_g XI10/NET3792
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2216 N_VSS_XI10/MM2216_d N_WL<55>_XI10/MM2216_g N_BL<12>_XI10/MM2216_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2252 N_VSS_XI10/MM2252_d N_WL<54>_XI10/MM2252_g XI10/NET4056
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2158 N_VSS_XI10/MM2158_d N_WL<53>_XI10/MM2158_g N_BL<12>_XI10/MM2158_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2134 N_VSS_XI10/MM2134_d N_WL<52>_XI10/MM2134_g XI10/NET3448
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2314 N_VSS_XI10/MM2314_d N_WL<51>_XI10/MM2314_g N_BL<12>_XI10/MM2314_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2290 N_VSS_XI10/MM2290_d N_WL<50>_XI10/MM2290_g XI10/NET3980
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2085 N_VSS_XI10/MM2085_d N_WL<49>_XI10/MM2085_g N_BL<12>_XI10/MM2085_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2116 N_VSS_XI10/MM2116_d N_WL<48>_XI10/MM2116_g XI10/NET3516
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2728 N_VSS_XI10/MM2728_d N_WL<47>_XI10/MM2728_g N_BL<12>_XI10/MM2728_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2764 N_VSS_XI10/MM2764_d N_WL<46>_XI10/MM2764_g XI10/NET4524
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2670 N_VSS_XI10/MM2670_d N_WL<45>_XI10/MM2670_g N_BL<12>_XI10/MM2670_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2646 N_VSS_XI10/MM2646_d N_WL<44>_XI10/MM2646_g XI10/NET4740
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2826 N_VSS_XI10/MM2826_d N_WL<43>_XI10/MM2826_g N_BL<12>_XI10/MM2826_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2802 N_VSS_XI10/MM2802_d N_WL<42>_XI10/MM2802_g XI10/NET4448
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2597 N_VSS_XI10/MM2597_d N_WL<41>_XI10/MM2597_g N_BL<12>_XI10/MM2597_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2694 N_VSS_XI10/MM2694_d N_WL<40>_XI10/MM2694_g XI10/NET4660
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2963 N_VSS_XI10/MM2963_d N_WL<39>_XI10/MM2963_g N_BL<12>_XI10/MM2963_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2938 N_VSS_XI10/MM2938_d N_WL<38>_XI10/MM2938_g XI10/NET5404
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3021 N_VSS_XI10/MM3021_d N_WL<37>_XI10/MM3021_g N_BL<12>_XI10/MM3021_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3056 N_VSS_XI10/MM3056_d N_WL<36>_XI10/MM3056_g XI10/NET5188
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2865 N_VSS_XI10/MM2865_d N_WL<35>_XI10/MM2865_g N_BL<12>_XI10/MM2865_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2900 N_VSS_XI10/MM2900_d N_WL<34>_XI10/MM2900_g XI10/NET4280
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3094 N_VSS_XI10/MM3094_d N_WL<33>_XI10/MM3094_g N_BL<12>_XI10/MM3094_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3063 N_VSS_XI10/MM3063_d N_WL<32>_XI10/MM3063_g XI10/NET5164
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1704 N_VSS_XI10/MM1704_d N_WL<31>_XI10/MM1704_g N_BL<12>_XI10/MM1704_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1740 N_VSS_XI10/MM1740_d N_WL<30>_XI10/MM1740_g XI10/NET2088
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1646 N_VSS_XI10/MM1646_d N_WL<29>_XI10/MM1646_g N_BL<12>_XI10/MM1646_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1622 N_VSS_XI10/MM1622_d N_WL<28>_XI10/MM1622_g XI10/NET2304
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1802 N_VSS_XI10/MM1802_d N_WL<27>_XI10/MM1802_g N_BL<12>_XI10/MM1802_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1778 N_VSS_XI10/MM1778_d N_WL<26>_XI10/MM1778_g XI10/NET2012
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1573 N_VSS_XI10/MM1573_d N_WL<25>_XI10/MM1573_g N_BL<12>_XI10/MM1573_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1670 N_VSS_XI10/MM1670_d N_WL<24>_XI10/MM1670_g XI10/NET2224
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1939 N_VSS_XI10/MM1939_d N_WL<23>_XI10/MM1939_g N_BL<12>_XI10/MM1939_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1914 N_VSS_XI10/MM1914_d N_WL<22>_XI10/MM1914_g XI10/NET2792
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1997 N_VSS_XI10/MM1997_d N_WL<21>_XI10/MM1997_g N_BL<12>_XI10/MM1997_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2032 N_VSS_XI10/MM2032_d N_WL<20>_XI10/MM2032_g XI10/NET02600
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1841 N_VSS_XI10/MM1841_d N_WL<19>_XI10/MM1841_g N_BL<12>_XI10/MM1841_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1876 N_VSS_XI10/MM1876_d N_WL<18>_XI10/MM1876_g XI10/NET2868
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2070 N_VSS_XI10/MM2070_d N_WL<17>_XI10/MM2070_g N_BL<12>_XI10/MM2070_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2061 N_VSS_XI10/MM2061_d N_WL<16>_XI10/MM2061_g XI10/NET2480
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1427 N_VSS_XI10/MM1427_d N_WL<15>_XI10/MM1427_g N_BL<12>_XI10/MM1427_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1391 N_VSS_XI10/MM1391_d N_WL<14>_XI10/MM1391_g XI10/NET5584
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1485 N_VSS_XI10/MM1485_d N_WL<13>_XI10/MM1485_g N_BL<12>_XI10/MM1485_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1520 N_VSS_XI10/MM1520_d N_WL<12>_XI10/MM1520_g XI10/NET1824
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1329 N_VSS_XI10/MM1329_d N_WL<11>_XI10/MM1329_g N_BL<12>_XI10/MM1329_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1353 N_VSS_XI10/MM1353_d N_WL<10>_XI10/MM1353_g XI10/NET5508
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1558 N_VSS_XI10/MM1558_d N_WL<9>_XI10/MM1558_g N_BL<12>_XI10/MM1558_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1549 N_VSS_XI10/MM1549_d N_WL<8>_XI10/MM1549_g XI10/NET1728
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1219 N_VSS_XI10/MM1219_d N_WL<7>_XI10/MM1219_g N_BL<12>_XI10/MM1219_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1184 N_VSS_XI10/MM1184_d N_WL<6>_XI10/MM1184_g XI10/NET3040
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1272 N_VSS_XI10/MM1272_d N_WL<5>_XI10/MM1272_g N_BL<12>_XI10/MM1272_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1296 N_VSS_XI10/MM1296_d N_WL<4>_XI10/MM1296_g XI10/NET3256
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1144 N_VSS_XI10/MM1144_d N_WL<3>_XI10/MM1144_g N_BL<12>_XI10/MM1144_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1168 N_VSS_XI10/MM1168_d N_WL<2>_XI10/MM1168_g XI10/NET1940
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1104 N_VSS_XI10/MM1104_d N_WL<1>_XI10/MM1104_g N_BL<12>_XI10/MM1104_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1067 N_VSS_XI10/MM1067_d N_WL<0>_XI10/MM1067_g XI10/NET3176
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI17/XI16/XI1/MM10 N_XI17/XI16/NET40_XI17/XI16/XI1/MM10_d
+ N_YOUT<5>_XI17/XI16/XI1/MM10_g N_VSS_XI17/XI16/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI15/XI1/MM10 N_XI17/XI15/NET40_XI17/XI15/XI1/MM10_d
+ N_YOUT<4>_XI17/XI15/XI1/MM10_g N_VSS_XI17/XI15/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI16/MM1 N_BL<13>_XI17/XI16/MM1_d N_XI17/XI16/NET40_XI17/XI16/MM1_g
+ N_DL<1>_XI17/XI16/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI15/MM1 N_BL<12>_XI17/XI15/MM1_d N_XI17/XI15/NET40_XI17/XI15/MM1_g
+ N_DL<1>_XI17/XI15/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2471 N_VSS_XI10/MM2471_d N_WL<63>_XI10/MM2471_g XI10/NET3668
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2425 N_VSS_XI10/MM2425_d N_WL<62>_XI10/MM2425_g N_BL<13>_XI10/MM2425_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2491 N_VSS_XI10/MM2491_d N_WL<61>_XI10/MM2491_g XI10/NET3624
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2534 N_VSS_XI10/MM2534_d N_WL<60>_XI10/MM2534_g N_BL<13>_XI10/MM2534_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2345 N_VSS_XI10/MM2345_d N_WL<59>_XI10/MM2345_g XI10/NET3876
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2378 N_VSS_XI10/MM2378_d N_WL<58>_XI10/MM2378_g N_BL<13>_XI10/MM2378_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2402 N_VSS_XI10/MM2402_d N_WL<57>_XI10/MM2402_g XI10/NET3800
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2490 N_VSS_XI10/MM2490_d N_WL<56>_XI10/MM2490_g N_BL<13>_XI10/MM2490_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2208 N_VSS_XI10/MM2208_d N_WL<55>_XI10/MM2208_g XI10/NET4124
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2242 N_VSS_XI10/MM2242_d N_WL<54>_XI10/MM2242_g N_BL<13>_XI10/MM2242_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2183 N_VSS_XI10/MM2183_d N_WL<53>_XI10/MM2183_g XI10/NET4188
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2133 N_VSS_XI10/MM2133_d N_WL<52>_XI10/MM2133_g N_BL<13>_XI10/MM2133_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2097 N_VSS_XI10/MM2097_d N_WL<51>_XI10/MM2097_g XI10/NET3584
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2289 N_VSS_XI10/MM2289_d N_WL<50>_XI10/MM2289_g N_BL<13>_XI10/MM2289_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2110 N_VSS_XI10/MM2110_d N_WL<49>_XI10/MM2110_g XI10/NET3540
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2177 N_VSS_XI10/MM2177_d N_WL<48>_XI10/MM2177_g N_BL<13>_XI10/MM2177_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2720 N_VSS_XI10/MM2720_d N_WL<47>_XI10/MM2720_g XI10/NET4592
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2754 N_VSS_XI10/MM2754_d N_WL<46>_XI10/MM2754_g N_BL<13>_XI10/MM2754_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2695 N_VSS_XI10/MM2695_d N_WL<45>_XI10/MM2695_g XI10/NET4656
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2645 N_VSS_XI10/MM2645_d N_WL<44>_XI10/MM2645_g N_BL<13>_XI10/MM2645_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2841 N_VSS_XI10/MM2841_d N_WL<43>_XI10/MM2841_g XI10/NET4400
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2801 N_VSS_XI10/MM2801_d N_WL<42>_XI10/MM2801_g N_BL<13>_XI10/MM2801_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2743 N_VSS_XI10/MM2743_d N_WL<41>_XI10/MM2743_g XI10/NET4580
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2689 N_VSS_XI10/MM2689_d N_WL<40>_XI10/MM2689_g N_BL<13>_XI10/MM2689_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2983 N_VSS_XI10/MM2983_d N_WL<39>_XI10/MM2983_g XI10/NET5336
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2937 N_VSS_XI10/MM2937_d N_WL<38>_XI10/MM2937_g N_BL<13>_XI10/MM2937_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3012 N_VSS_XI10/MM3012_d N_WL<37>_XI10/MM3012_g XI10/NET5256
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3046 N_VSS_XI10/MM3046_d N_WL<36>_XI10/MM3046_g N_BL<13>_XI10/MM3046_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2857 N_VSS_XI10/MM2857_d N_WL<35>_XI10/MM2857_g XI10/NET4344
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2890 N_VSS_XI10/MM2890_d N_WL<34>_XI10/MM2890_g N_BL<13>_XI10/MM2890_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3077 N_VSS_XI10/MM3077_d N_WL<33>_XI10/MM3077_g XI10/NET5108
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3002 N_VSS_XI10/MM3002_d N_WL<32>_XI10/MM3002_g N_BL<13>_XI10/MM3002_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1696 N_VSS_XI10/MM1696_d N_WL<31>_XI10/MM1696_g XI10/NET2156
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1730 N_VSS_XI10/MM1730_d N_WL<30>_XI10/MM1730_g N_BL<13>_XI10/MM1730_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1671 N_VSS_XI10/MM1671_d N_WL<29>_XI10/MM1671_g XI10/NET2220
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1621 N_VSS_XI10/MM1621_d N_WL<28>_XI10/MM1621_g N_BL<13>_XI10/MM1621_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1591 N_VSS_XI10/MM1591_d N_WL<27>_XI10/MM1591_g XI10/NET2424
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1777 N_VSS_XI10/MM1777_d N_WL<26>_XI10/MM1777_g N_BL<13>_XI10/MM1777_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1719 N_VSS_XI10/MM1719_d N_WL<25>_XI10/MM1719_g XI10/NET2144
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1665 N_VSS_XI10/MM1665_d N_WL<24>_XI10/MM1665_g N_BL<13>_XI10/MM1665_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1959 N_VSS_XI10/MM1959_d N_WL<23>_XI10/MM1959_g XI10/NET2724
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1913 N_VSS_XI10/MM1913_d N_WL<22>_XI10/MM1913_g N_BL<13>_XI10/MM1913_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1988 N_VSS_XI10/MM1988_d N_WL<21>_XI10/MM1988_g XI10/NET2644
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2022 N_VSS_XI10/MM2022_d N_WL<20>_XI10/MM2022_g N_BL<13>_XI10/MM2022_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2052 N_VSS_XI10/MM2052_d N_WL<19>_XI10/MM2052_g XI10/NET2500
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1866 N_VSS_XI10/MM1866_d N_WL<18>_XI10/MM1866_g N_BL<13>_XI10/MM1866_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2053 N_VSS_XI10/MM2053_d N_WL<17>_XI10/MM2053_g XI10/NET2496
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1978 N_VSS_XI10/MM1978_d N_WL<16>_XI10/MM1978_g N_BL<13>_XI10/MM1978_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1435 N_VSS_XI10/MM1435_d N_WL<15>_XI10/MM1435_g XI10/NET5652
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1401 N_VSS_XI10/MM1401_d N_WL<14>_XI10/MM1401_g N_BL<13>_XI10/MM1401_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1460 N_VSS_XI10/MM1460_d N_WL<13>_XI10/MM1460_g XI10/NET5720
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1510 N_VSS_XI10/MM1510_d N_WL<12>_XI10/MM1510_g N_BL<13>_XI10/MM1510_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1540 N_VSS_XI10/MM1540_d N_WL<11>_XI10/MM1540_g XI10/NET1748
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1354 N_VSS_XI10/MM1354_d N_WL<10>_XI10/MM1354_g N_BL<13>_XI10/MM1354_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1541 N_VSS_XI10/MM1541_d N_WL<9>_XI10/MM1541_g XI10/NET1744
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1466 N_VSS_XI10/MM1466_d N_WL<8>_XI10/MM1466_g N_BL<13>_XI10/MM1466_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1227 N_VSS_XI10/MM1227_d N_WL<7>_XI10/MM1227_g XI10/NET3108
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1194 N_VSS_XI10/MM1194_d N_WL<6>_XI10/MM1194_g N_BL<13>_XI10/MM1194_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1252 N_VSS_XI10/MM1252_d N_WL<5>_XI10/MM1252_g XI10/NET3172
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1297 N_VSS_XI10/MM1297_d N_WL<4>_XI10/MM1297_g N_BL<13>_XI10/MM1297_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1129 N_VSS_XI10/MM1129_d N_WL<3>_XI10/MM1129_g XI10/NET1892
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1169 N_VSS_XI10/MM1169_d N_WL<2>_XI10/MM1169_g N_BL<13>_XI10/MM1169_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1105 N_VSS_XI10/MM1105_d N_WL<1>_XI10/MM1105_g XI10/NET3096
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1066 N_VSS_XI10/MM1066_d N_WL<0>_XI10/MM1066_g N_BL<13>_XI10/MM1066_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2476 N_VSS_XI10/MM2476_d N_WL<63>_XI10/MM2476_g N_BL<14>_XI10/MM2476_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2413 N_VSS_XI10/MM2413_d N_WL<62>_XI10/MM2413_g XI10/NET3788
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2479 N_VSS_XI10/MM2479_d N_WL<61>_XI10/MM2479_g N_BL<14>_XI10/MM2479_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2546 N_VSS_XI10/MM2546_d N_WL<60>_XI10/MM2546_g XI10/NET5004
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2508 N_VSS_XI10/MM2508_d N_WL<59>_XI10/MM2508_g N_BL<14>_XI10/MM2508_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2390 N_VSS_XI10/MM2390_d N_WL<58>_XI10/MM2390_g XI10/NET3804
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2335 N_VSS_XI10/MM2335_d N_WL<57>_XI10/MM2335_g N_BL<14>_XI10/MM2335_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2485 N_VSS_XI10/MM2485_d N_WL<56>_XI10/MM2485_g XI10/NET3644
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2191 N_VSS_XI10/MM2191_d N_WL<55>_XI10/MM2191_g N_BL<14>_XI10/MM2191_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2254 N_VSS_XI10/MM2254_d N_WL<54>_XI10/MM2254_g XI10/NET4048
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2188 N_VSS_XI10/MM2188_d N_WL<53>_XI10/MM2188_g N_BL<14>_XI10/MM2188_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2135 N_VSS_XI10/MM2135_d N_WL<52>_XI10/MM2135_g XI10/NET3444
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2159 N_VSS_XI10/MM2159_d N_WL<51>_XI10/MM2159_g N_BL<14>_XI10/MM2159_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2291 N_VSS_XI10/MM2291_d N_WL<50>_XI10/MM2291_g XI10/NET3976
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2332 N_VSS_XI10/MM2332_d N_WL<49>_XI10/MM2332_g N_BL<14>_XI10/MM2332_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2120 N_VSS_XI10/MM2120_d N_WL<48>_XI10/MM2120_g XI10/NET3504
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2703 N_VSS_XI10/MM2703_d N_WL<47>_XI10/MM2703_g N_BL<14>_XI10/MM2703_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2766 N_VSS_XI10/MM2766_d N_WL<46>_XI10/MM2766_g XI10/NET4516
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2700 N_VSS_XI10/MM2700_d N_WL<45>_XI10/MM2700_g N_BL<14>_XI10/MM2700_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2647 N_VSS_XI10/MM2647_d N_WL<44>_XI10/MM2647_g XI10/NET4736
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2671 N_VSS_XI10/MM2671_d N_WL<43>_XI10/MM2671_g N_BL<14>_XI10/MM2671_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2803 N_VSS_XI10/MM2803_d N_WL<42>_XI10/MM2803_g XI10/NET4444
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2844 N_VSS_XI10/MM2844_d N_WL<41>_XI10/MM2844_g N_BL<14>_XI10/MM2844_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2767 N_VSS_XI10/MM2767_d N_WL<40>_XI10/MM2767_g XI10/NET4512
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2988 N_VSS_XI10/MM2988_d N_WL<39>_XI10/MM2988_g N_BL<14>_XI10/MM2988_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2939 N_VSS_XI10/MM2939_d N_WL<38>_XI10/MM2939_g XI10/NET5400
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2991 N_VSS_XI10/MM2991_d N_WL<37>_XI10/MM2991_g N_BL<14>_XI10/MM2991_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3058 N_VSS_XI10/MM3058_d N_WL<36>_XI10/MM3058_g XI10/NET5180
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3020 N_VSS_XI10/MM3020_d N_WL<35>_XI10/MM3020_g N_BL<14>_XI10/MM3020_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2902 N_VSS_XI10/MM2902_d N_WL<34>_XI10/MM2902_g XI10/NET4272
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2847 N_VSS_XI10/MM2847_d N_WL<33>_XI10/MM2847_g N_BL<14>_XI10/MM2847_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3064 N_VSS_XI10/MM3064_d N_WL<32>_XI10/MM3064_g XI10/NET5160
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1679 N_VSS_XI10/MM1679_d N_WL<31>_XI10/MM1679_g N_BL<14>_XI10/MM1679_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1742 N_VSS_XI10/MM1742_d N_WL<30>_XI10/MM1742_g XI10/NET2080
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1676 N_VSS_XI10/MM1676_d N_WL<29>_XI10/MM1676_g N_BL<14>_XI10/MM1676_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1623 N_VSS_XI10/MM1623_d N_WL<28>_XI10/MM1623_g XI10/NET2300
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1647 N_VSS_XI10/MM1647_d N_WL<27>_XI10/MM1647_g N_BL<14>_XI10/MM1647_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1779 N_VSS_XI10/MM1779_d N_WL<26>_XI10/MM1779_g XI10/NET2008
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1820 N_VSS_XI10/MM1820_d N_WL<25>_XI10/MM1820_g N_BL<14>_XI10/MM1820_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1743 N_VSS_XI10/MM1743_d N_WL<24>_XI10/MM1743_g XI10/NET2076
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1964 N_VSS_XI10/MM1964_d N_WL<23>_XI10/MM1964_g N_BL<14>_XI10/MM1964_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1915 N_VSS_XI10/MM1915_d N_WL<22>_XI10/MM1915_g XI10/NET2788
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1967 N_VSS_XI10/MM1967_d N_WL<21>_XI10/MM1967_g N_BL<14>_XI10/MM1967_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2034 N_VSS_XI10/MM2034_d N_WL<20>_XI10/MM2034_g XI10/NET02592
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1996 N_VSS_XI10/MM1996_d N_WL<19>_XI10/MM1996_g N_BL<14>_XI10/MM1996_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1878 N_VSS_XI10/MM1878_d N_WL<18>_XI10/MM1878_g XI10/NET2860
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1823 N_VSS_XI10/MM1823_d N_WL<17>_XI10/MM1823_g N_BL<14>_XI10/MM1823_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2077 N_VSS_XI10/MM2077_d N_WL<16>_XI10/MM2077_g XI10/NET2464
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1452 N_VSS_XI10/MM1452_d N_WL<15>_XI10/MM1452_g N_BL<14>_XI10/MM1452_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1389 N_VSS_XI10/MM1389_d N_WL<14>_XI10/MM1389_g XI10/NET5576
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1455 N_VSS_XI10/MM1455_d N_WL<13>_XI10/MM1455_g N_BL<14>_XI10/MM1455_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1522 N_VSS_XI10/MM1522_d N_WL<12>_XI10/MM1522_g XI10/NET1816
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1484 N_VSS_XI10/MM1484_d N_WL<11>_XI10/MM1484_g N_BL<14>_XI10/MM1484_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1352 N_VSS_XI10/MM1352_d N_WL<10>_XI10/MM1352_g XI10/NET5504
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1311 N_VSS_XI10/MM1311_d N_WL<9>_XI10/MM1311_g N_BL<14>_XI10/MM1311_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1565 N_VSS_XI10/MM1565_d N_WL<8>_XI10/MM1565_g XI10/NET1712
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1244 N_VSS_XI10/MM1244_d N_WL<7>_XI10/MM1244_g N_BL<14>_XI10/MM1244_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1182 N_VSS_XI10/MM1182_d N_WL<6>_XI10/MM1182_g XI10/NET3032
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1247 N_VSS_XI10/MM1247_d N_WL<5>_XI10/MM1247_g N_BL<14>_XI10/MM1247_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1295 N_VSS_XI10/MM1295_d N_WL<4>_XI10/MM1295_g XI10/NET3252
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1119 N_VSS_XI10/MM1119_d N_WL<3>_XI10/MM1119_g N_BL<14>_XI10/MM1119_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1167 N_VSS_XI10/MM1167_d N_WL<2>_XI10/MM1167_g XI10/NET1936
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1103 N_VSS_XI10/MM1103_d N_WL<1>_XI10/MM1103_g N_BL<14>_XI10/MM1103_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1068 N_VSS_XI10/MM1068_d N_WL<0>_XI10/MM1068_g XI10/NET3028
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI17/XI18/XI1/MM10 N_XI17/XI18/NET40_XI17/XI18/XI1/MM10_d
+ N_YOUT<7>_XI17/XI18/XI1/MM10_g N_VSS_XI17/XI18/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI17/XI1/MM10 N_XI17/XI17/NET40_XI17/XI17/XI1/MM10_d
+ N_YOUT<6>_XI17/XI17/XI1/MM10_g N_VSS_XI17/XI17/XI1/MM10_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI18/MM1 N_BL<15>_XI17/XI18/MM1_d N_XI17/XI18/NET40_XI17/XI18/MM1_g
+ N_DL<1>_XI17/XI18/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI17/XI17/MM1 N_BL<14>_XI17/XI17/MM1_d N_XI17/XI17/NET40_XI17/XI17/MM1_g
+ N_DL<1>_XI17/XI17/MM1_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI10/MM2472 N_VSS_XI10/MM2472_d N_WL<63>_XI10/MM2472_g XI10/NET3664
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2428 N_VSS_XI10/MM2428_d N_WL<62>_XI10/MM2428_g N_BL<15>_XI10/MM2428_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2495 N_VSS_XI10/MM2495_d N_WL<61>_XI10/MM2495_g XI10/NET3608
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2531 N_VSS_XI10/MM2531_d N_WL<60>_XI10/MM2531_g N_BL<15>_XI10/MM2531_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2357 N_VSS_XI10/MM2357_d N_WL<59>_XI10/MM2357_g XI10/NET3868
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2375 N_VSS_XI10/MM2375_d N_WL<58>_XI10/MM2375_g N_BL<15>_XI10/MM2375_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2436 N_VSS_XI10/MM2436_d N_WL<57>_XI10/MM2436_g XI10/NET3724
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2411 N_VSS_XI10/MM2411_d N_WL<56>_XI10/MM2411_g N_BL<15>_XI10/MM2411_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2220 N_VSS_XI10/MM2220_d N_WL<55>_XI10/MM2220_g XI10/NET4116
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2239 N_VSS_XI10/MM2239_d N_WL<54>_XI10/MM2239_g N_BL<15>_XI10/MM2239_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2184 N_VSS_XI10/MM2184_d N_WL<53>_XI10/MM2184_g XI10/NET4184
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2136 N_VSS_XI10/MM2136_d N_WL<52>_XI10/MM2136_g N_BL<15>_XI10/MM2136_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2103 N_VSS_XI10/MM2103_d N_WL<51>_XI10/MM2103_g XI10/NET3568
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2292 N_VSS_XI10/MM2292_d N_WL<50>_XI10/MM2292_g N_BL<15>_XI10/MM2292_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2111 N_VSS_XI10/MM2111_d N_WL<49>_XI10/MM2111_g XI10/NET3536
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2256 N_VSS_XI10/MM2256_d N_WL<48>_XI10/MM2256_g N_BL<15>_XI10/MM2256_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2732 N_VSS_XI10/MM2732_d N_WL<47>_XI10/MM2732_g XI10/NET4584
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2751 N_VSS_XI10/MM2751_d N_WL<46>_XI10/MM2751_g N_BL<15>_XI10/MM2751_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2696 N_VSS_XI10/MM2696_d N_WL<45>_XI10/MM2696_g XI10/NET4652
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2648 N_VSS_XI10/MM2648_d N_WL<44>_XI10/MM2648_g N_BL<15>_XI10/MM2648_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2842 N_VSS_XI10/MM2842_d N_WL<43>_XI10/MM2842_g XI10/NET4396
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2804 N_VSS_XI10/MM2804_d N_WL<42>_XI10/MM2804_g N_BL<15>_XI10/MM2804_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2777 N_VSS_XI10/MM2777_d N_WL<41>_XI10/MM2777_g XI10/NET4504
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2768 N_VSS_XI10/MM2768_d N_WL<40>_XI10/MM2768_g N_BL<15>_XI10/MM2768_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2984 N_VSS_XI10/MM2984_d N_WL<39>_XI10/MM2984_g XI10/NET5332
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2940 N_VSS_XI10/MM2940_d N_WL<38>_XI10/MM2940_g N_BL<15>_XI10/MM2940_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3025 N_VSS_XI10/MM3025_d N_WL<37>_XI10/MM3025_g XI10/NET5244
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM3043 N_VSS_XI10/MM3043_d N_WL<36>_XI10/MM3043_g N_BL<15>_XI10/MM3043_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2869 N_VSS_XI10/MM2869_d N_WL<35>_XI10/MM2869_g XI10/NET4336
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2887 N_VSS_XI10/MM2887_d N_WL<34>_XI10/MM2887_g N_BL<15>_XI10/MM2887_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2914 N_VSS_XI10/MM2914_d N_WL<33>_XI10/MM2914_g XI10/NET4268
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2923 N_VSS_XI10/MM2923_d N_WL<32>_XI10/MM2923_g N_BL<15>_XI10/MM2923_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1708 N_VSS_XI10/MM1708_d N_WL<31>_XI10/MM1708_g XI10/NET2148
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1727 N_VSS_XI10/MM1727_d N_WL<30>_XI10/MM1727_g N_BL<15>_XI10/MM1727_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1672 N_VSS_XI10/MM1672_d N_WL<29>_XI10/MM1672_g XI10/NET2216
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1624 N_VSS_XI10/MM1624_d N_WL<28>_XI10/MM1624_g N_BL<15>_XI10/MM1624_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1798 N_VSS_XI10/MM1798_d N_WL<27>_XI10/MM1798_g XI10/NET2000
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1780 N_VSS_XI10/MM1780_d N_WL<26>_XI10/MM1780_g N_BL<15>_XI10/MM1780_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1753 N_VSS_XI10/MM1753_d N_WL<25>_XI10/MM1753_g XI10/NET2068
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1744 N_VSS_XI10/MM1744_d N_WL<24>_XI10/MM1744_g N_BL<15>_XI10/MM1744_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1960 N_VSS_XI10/MM1960_d N_WL<23>_XI10/MM1960_g XI10/NET2720
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1916 N_VSS_XI10/MM1916_d N_WL<22>_XI10/MM1916_g N_BL<15>_XI10/MM1916_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2001 N_VSS_XI10/MM2001_d N_WL<21>_XI10/MM2001_g XI10/NET2632
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2019 N_VSS_XI10/MM2019_d N_WL<20>_XI10/MM2019_g N_BL<15>_XI10/MM2019_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2058 N_VSS_XI10/MM2058_d N_WL<19>_XI10/MM2058_g XI10/NET2484
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1863 N_VSS_XI10/MM1863_d N_WL<18>_XI10/MM1863_g N_BL<15>_XI10/MM1863_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM2074 N_VSS_XI10/MM2074_d N_WL<17>_XI10/MM2074_g XI10/NET2472
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1899 N_VSS_XI10/MM1899_d N_WL<16>_XI10/MM1899_g N_BL<15>_XI10/MM1899_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1423 N_VSS_XI10/MM1423_d N_WL<15>_XI10/MM1423_g XI10/NET5644
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1404 N_VSS_XI10/MM1404_d N_WL<14>_XI10/MM1404_g N_BL<15>_XI10/MM1404_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1459 N_VSS_XI10/MM1459_d N_WL<13>_XI10/MM1459_g XI10/NET5716
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1507 N_VSS_XI10/MM1507_d N_WL<12>_XI10/MM1507_g N_BL<15>_XI10/MM1507_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1546 N_VSS_XI10/MM1546_d N_WL<11>_XI10/MM1546_g XI10/NET1732
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1351 N_VSS_XI10/MM1351_d N_WL<10>_XI10/MM1351_g N_BL<15>_XI10/MM1351_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1562 N_VSS_XI10/MM1562_d N_WL<9>_XI10/MM1562_g XI10/NET1720
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1387 N_VSS_XI10/MM1387_d N_WL<8>_XI10/MM1387_g N_BL<15>_XI10/MM1387_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1215 N_VSS_XI10/MM1215_d N_WL<7>_XI10/MM1215_g XI10/NET3100
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1197 N_VSS_XI10/MM1197_d N_WL<6>_XI10/MM1197_g N_BL<15>_XI10/MM1197_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1251 N_VSS_XI10/MM1251_d N_WL<5>_XI10/MM1251_g XI10/NET3168
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1294 N_VSS_XI10/MM1294_d N_WL<4>_XI10/MM1294_g N_BL<15>_XI10/MM1294_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1128 N_VSS_XI10/MM1128_d N_WL<3>_XI10/MM1128_g XI10/NET1888
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1166 N_VSS_XI10/MM1166_d N_WL<2>_XI10/MM1166_g N_BL<15>_XI10/MM1166_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1106 N_VSS_XI10/MM1106_d N_WL<1>_XI10/MM1106_g XI10/NET1996
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI10/MM1069 N_VSS_XI10/MM1069_d N_WL<0>_XI10/MM1069_g N_BL<15>_XI10/MM1069_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXI9/XI0/XI10/MM6 N_XI9/XI0/NET0116_XI9/XI0/XI10/MM6_d
+ N_X_SEL<3>_XI9/XI0/XI10/MM6_g N_VDD_XI9/XI0/XI10/MM6_s
+ N_VDD_XI9/XI0/XI10/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI9/XI0/XI11/MM6 N_XI9/XI0/NET0105_XI9/XI0/XI11/MM6_d
+ N_X_SEL<4>_XI9/XI0/XI11/MM6_g N_VDD_XI9/XI0/XI11/MM6_s
+ N_VDD_XI9/XI0/XI11/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI9/XI0/XI8/MM6 N_XI9/XI0/NET0158_XI9/XI0/XI8/MM6_d
+ N_X_SEL<5>_XI9/XI0/XI8/MM6_g N_VDD_XI9/XI0/XI8/MM6_s N_VDD_XI9/XI0/XI8/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI9/XI1/XI10/MM6 N_XI9/XI1/NET0116_XI9/XI1/XI10/MM6_d
+ N_X_SEL<0>_XI9/XI1/XI10/MM6_g N_VDD_XI9/XI1/XI10/MM6_s
+ N_VDD_XI9/XI1/XI10/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI9/XI1/XI11/MM6 N_XI9/XI1/NET0105_XI9/XI1/XI11/MM6_d
+ N_X_SEL<1>_XI9/XI1/XI11/MM6_g N_VDD_XI9/XI1/XI11/MM6_s
+ N_VDD_XI9/XI1/XI11/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI9/XI1/XI8/MM6 N_XI9/XI1/NET0158_XI9/XI1/XI8/MM6_d
+ N_X_SEL<2>_XI9/XI1/XI8/MM6_g N_VDD_XI9/XI1/XI8/MM6_s N_VDD_XI9/XI1/XI8/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI9/XI0/XI7/MM12 N_XI9/NET17_XI9/XI0/XI7/MM12_d N_WLEN_XI9/XI0/XI7/MM12_g
+ N_VDD_XI9/XI0/XI7/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI7/MM2 N_XI9/NET17_XI9/XI0/XI7/MM2_d N_X_SEL<3>_XI9/XI0/XI7/MM2_g
+ N_VDD_XI9/XI0/XI7/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI7/MM0 N_XI9/NET17_XI9/XI0/XI7/MM0_d N_X_SEL<4>_XI9/XI0/XI7/MM0_g
+ N_VDD_XI9/XI0/XI7/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI7/MM10 N_XI9/NET17_XI9/XI0/XI7/MM10_d N_X_SEL<5>_XI9/XI0/XI7/MM10_g
+ N_VDD_XI9/XI0/XI7/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI6/MM12 N_XI9/NET18_XI9/XI0/XI6/MM12_d N_WLEN_XI9/XI0/XI6/MM12_g
+ N_VDD_XI9/XI0/XI6/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI6/MM2 N_XI9/NET18_XI9/XI0/XI6/MM2_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI6/MM2_g N_VDD_XI9/XI0/XI6/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI6/MM0 N_XI9/NET18_XI9/XI0/XI6/MM0_d N_X_SEL<4>_XI9/XI0/XI6/MM0_g
+ N_VDD_XI9/XI0/XI6/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI6/MM10 N_XI9/NET18_XI9/XI0/XI6/MM10_d N_X_SEL<5>_XI9/XI0/XI6/MM10_g
+ N_VDD_XI9/XI0/XI6/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI5/MM12 N_XI9/NET19_XI9/XI0/XI5/MM12_d N_WLEN_XI9/XI0/XI5/MM12_g
+ N_VDD_XI9/XI0/XI5/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI5/MM2 N_XI9/NET19_XI9/XI0/XI5/MM2_d N_X_SEL<3>_XI9/XI0/XI5/MM2_g
+ N_VDD_XI9/XI0/XI5/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI5/MM0 N_XI9/NET19_XI9/XI0/XI5/MM0_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI5/MM0_g N_VDD_XI9/XI0/XI5/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI5/MM10 N_XI9/NET19_XI9/XI0/XI5/MM10_d N_X_SEL<5>_XI9/XI0/XI5/MM10_g
+ N_VDD_XI9/XI0/XI5/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI4/MM12 N_XI9/NET20_XI9/XI0/XI4/MM12_d N_WLEN_XI9/XI0/XI4/MM12_g
+ N_VDD_XI9/XI0/XI4/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI4/MM2 N_XI9/NET20_XI9/XI0/XI4/MM2_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI4/MM2_g N_VDD_XI9/XI0/XI4/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI4/MM0 N_XI9/NET20_XI9/XI0/XI4/MM0_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI4/MM0_g N_VDD_XI9/XI0/XI4/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI4/MM10 N_XI9/NET20_XI9/XI0/XI4/MM10_d N_X_SEL<5>_XI9/XI0/XI4/MM10_g
+ N_VDD_XI9/XI0/XI4/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI3/MM12 N_XI9/NET21_XI9/XI0/XI3/MM12_d N_WLEN_XI9/XI0/XI3/MM12_g
+ N_VDD_XI9/XI0/XI3/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI3/MM2 N_XI9/NET21_XI9/XI0/XI3/MM2_d N_X_SEL<3>_XI9/XI0/XI3/MM2_g
+ N_VDD_XI9/XI0/XI3/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI3/MM0 N_XI9/NET21_XI9/XI0/XI3/MM0_d N_X_SEL<4>_XI9/XI0/XI3/MM0_g
+ N_VDD_XI9/XI0/XI3/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI3/MM10 N_XI9/NET21_XI9/XI0/XI3/MM10_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI3/MM10_g N_VDD_XI9/XI0/XI3/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI2/MM12 N_XI9/NET22_XI9/XI0/XI2/MM12_d N_WLEN_XI9/XI0/XI2/MM12_g
+ N_VDD_XI9/XI0/XI2/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI2/MM2 N_XI9/NET22_XI9/XI0/XI2/MM2_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI2/MM2_g N_VDD_XI9/XI0/XI2/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI2/MM0 N_XI9/NET22_XI9/XI0/XI2/MM0_d N_X_SEL<4>_XI9/XI0/XI2/MM0_g
+ N_VDD_XI9/XI0/XI2/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI2/MM10 N_XI9/NET22_XI9/XI0/XI2/MM10_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI2/MM10_g N_VDD_XI9/XI0/XI2/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI1/MM12 N_XI9/NET23_XI9/XI0/XI1/MM12_d N_WLEN_XI9/XI0/XI1/MM12_g
+ N_VDD_XI9/XI0/XI1/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI1/MM2 N_XI9/NET23_XI9/XI0/XI1/MM2_d N_X_SEL<3>_XI9/XI0/XI1/MM2_g
+ N_VDD_XI9/XI0/XI1/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI1/MM0 N_XI9/NET23_XI9/XI0/XI1/MM0_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI1/MM0_g N_VDD_XI9/XI0/XI1/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI1/MM10 N_XI9/NET23_XI9/XI0/XI1/MM10_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI1/MM10_g N_VDD_XI9/XI0/XI1/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI0/MM12 N_XI9/NET24_XI9/XI0/XI0/MM12_d N_WLEN_XI9/XI0/XI0/MM12_g
+ N_VDD_XI9/XI0/XI0/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI0/MM2 N_XI9/NET24_XI9/XI0/XI0/MM2_d
+ N_XI9/XI0/NET0116_XI9/XI0/XI0/MM2_g N_VDD_XI9/XI0/XI0/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI0/MM0 N_XI9/NET24_XI9/XI0/XI0/MM0_d
+ N_XI9/XI0/NET0105_XI9/XI0/XI0/MM0_g N_VDD_XI9/XI0/XI0/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI0/XI0/MM10 N_XI9/NET24_XI9/XI0/XI0/MM10_d
+ N_XI9/XI0/NET0158_XI9/XI0/XI0/MM10_g N_VDD_XI9/XI0/XI0/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI7/MM12 N_XI9/NET4_XI9/XI1/XI7/MM12_d N_WLEN_XI9/XI1/XI7/MM12_g
+ N_VDD_XI9/XI1/XI7/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI7/MM2 N_XI9/NET4_XI9/XI1/XI7/MM2_d N_X_SEL<0>_XI9/XI1/XI7/MM2_g
+ N_VDD_XI9/XI1/XI7/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI7/MM0 N_XI9/NET4_XI9/XI1/XI7/MM0_d N_X_SEL<1>_XI9/XI1/XI7/MM0_g
+ N_VDD_XI9/XI1/XI7/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI7/MM10 N_XI9/NET4_XI9/XI1/XI7/MM10_d N_X_SEL<2>_XI9/XI1/XI7/MM10_g
+ N_VDD_XI9/XI1/XI7/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI6/MM12 N_XI9/NET5_XI9/XI1/XI6/MM12_d N_WLEN_XI9/XI1/XI6/MM12_g
+ N_VDD_XI9/XI1/XI6/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI6/MM2 N_XI9/NET5_XI9/XI1/XI6/MM2_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI6/MM2_g N_VDD_XI9/XI1/XI6/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI6/MM0 N_XI9/NET5_XI9/XI1/XI6/MM0_d N_X_SEL<1>_XI9/XI1/XI6/MM0_g
+ N_VDD_XI9/XI1/XI6/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI6/MM10 N_XI9/NET5_XI9/XI1/XI6/MM10_d N_X_SEL<2>_XI9/XI1/XI6/MM10_g
+ N_VDD_XI9/XI1/XI6/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI5/MM12 N_XI9/NET6_XI9/XI1/XI5/MM12_d N_WLEN_XI9/XI1/XI5/MM12_g
+ N_VDD_XI9/XI1/XI5/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI5/MM2 N_XI9/NET6_XI9/XI1/XI5/MM2_d N_X_SEL<0>_XI9/XI1/XI5/MM2_g
+ N_VDD_XI9/XI1/XI5/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI5/MM0 N_XI9/NET6_XI9/XI1/XI5/MM0_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI5/MM0_g N_VDD_XI9/XI1/XI5/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI5/MM10 N_XI9/NET6_XI9/XI1/XI5/MM10_d N_X_SEL<2>_XI9/XI1/XI5/MM10_g
+ N_VDD_XI9/XI1/XI5/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI4/MM12 N_XI9/NET7_XI9/XI1/XI4/MM12_d N_WLEN_XI9/XI1/XI4/MM12_g
+ N_VDD_XI9/XI1/XI4/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI4/MM2 N_XI9/NET7_XI9/XI1/XI4/MM2_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI4/MM2_g N_VDD_XI9/XI1/XI4/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI4/MM0 N_XI9/NET7_XI9/XI1/XI4/MM0_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI4/MM0_g N_VDD_XI9/XI1/XI4/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI4/MM10 N_XI9/NET7_XI9/XI1/XI4/MM10_d N_X_SEL<2>_XI9/XI1/XI4/MM10_g
+ N_VDD_XI9/XI1/XI4/MM10_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI3/MM12 N_XI9/NET8_XI9/XI1/XI3/MM12_d N_WLEN_XI9/XI1/XI3/MM12_g
+ N_VDD_XI9/XI1/XI3/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI3/MM2 N_XI9/NET8_XI9/XI1/XI3/MM2_d N_X_SEL<0>_XI9/XI1/XI3/MM2_g
+ N_VDD_XI9/XI1/XI3/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI3/MM0 N_XI9/NET8_XI9/XI1/XI3/MM0_d N_X_SEL<1>_XI9/XI1/XI3/MM0_g
+ N_VDD_XI9/XI1/XI3/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI3/MM10 N_XI9/NET8_XI9/XI1/XI3/MM10_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI3/MM10_g N_VDD_XI9/XI1/XI3/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI2/MM12 N_XI9/NET9_XI9/XI1/XI2/MM12_d N_WLEN_XI9/XI1/XI2/MM12_g
+ N_VDD_XI9/XI1/XI2/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI2/MM2 N_XI9/NET9_XI9/XI1/XI2/MM2_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI2/MM2_g N_VDD_XI9/XI1/XI2/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI2/MM0 N_XI9/NET9_XI9/XI1/XI2/MM0_d N_X_SEL<1>_XI9/XI1/XI2/MM0_g
+ N_VDD_XI9/XI1/XI2/MM0_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI2/MM10 N_XI9/NET9_XI9/XI1/XI2/MM10_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI2/MM10_g N_VDD_XI9/XI1/XI2/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI1/MM12 N_XI9/NET10_XI9/XI1/XI1/MM12_d N_WLEN_XI9/XI1/XI1/MM12_g
+ N_VDD_XI9/XI1/XI1/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI1/MM2 N_XI9/NET10_XI9/XI1/XI1/MM2_d N_X_SEL<0>_XI9/XI1/XI1/MM2_g
+ N_VDD_XI9/XI1/XI1/MM2_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI1/MM0 N_XI9/NET10_XI9/XI1/XI1/MM0_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI1/MM0_g N_VDD_XI9/XI1/XI1/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI1/MM10 N_XI9/NET10_XI9/XI1/XI1/MM10_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI1/MM10_g N_VDD_XI9/XI1/XI1/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI0/MM12 N_XI9/NET11_XI9/XI1/XI0/MM12_d N_WLEN_XI9/XI1/XI0/MM12_g
+ N_VDD_XI9/XI1/XI0/MM12_s N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI0/MM2 N_XI9/NET11_XI9/XI1/XI0/MM2_d
+ N_XI9/XI1/NET0116_XI9/XI1/XI0/MM2_g N_VDD_XI9/XI1/XI0/MM2_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI0/MM0 N_XI9/NET11_XI9/XI1/XI0/MM0_d
+ N_XI9/XI1/NET0105_XI9/XI1/XI0/MM0_g N_VDD_XI9/XI1/XI0/MM0_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI1/XI0/MM10 N_XI9/NET11_XI9/XI1/XI0/MM10_d
+ N_XI9/XI1/NET0158_XI9/XI1/XI0/MM10_g N_VDD_XI9/XI1/XI0/MM10_s
+ N_VDD_XI9/XI0/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9/XI136/MM0 N_WL<63>_XI9/XI136/MM0_d N_XI9/NET17_XI9/XI136/MM0_g
+ N_XI9/XI136/NET043_XI9/XI136/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI135/MM0 N_WL<62>_XI9/XI135/MM0_d N_XI9/NET17_XI9/XI135/MM0_g
+ N_XI9/XI135/NET043_XI9/XI135/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI137/MM0 N_WL<61>_XI9/XI137/MM0_d N_XI9/NET17_XI9/XI137/MM0_g
+ N_XI9/XI137/NET043_XI9/XI137/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI138/MM0 N_WL<60>_XI9/XI138/MM0_d N_XI9/NET17_XI9/XI138/MM0_g
+ N_XI9/XI138/NET043_XI9/XI138/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI133/MM0 N_WL<59>_XI9/XI133/MM0_d N_XI9/NET17_XI9/XI133/MM0_g
+ N_XI9/XI133/NET043_XI9/XI133/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI134/MM0 N_WL<58>_XI9/XI134/MM0_d N_XI9/NET17_XI9/XI134/MM0_g
+ N_XI9/XI134/NET043_XI9/XI134/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI132/MM0 N_WL<57>_XI9/XI132/MM0_d N_XI9/NET17_XI9/XI132/MM0_g
+ N_XI9/XI132/NET043_XI9/XI132/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI131/MM0 N_WL<56>_XI9/XI131/MM0_d N_XI9/NET17_XI9/XI131/MM0_g
+ N_XI9/XI131/NET043_XI9/XI131/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI141/MM0 N_WL<55>_XI9/XI141/MM0_d N_XI9/NET18_XI9/XI141/MM0_g
+ N_XI9/XI141/NET043_XI9/XI141/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI142/MM0 N_WL<54>_XI9/XI142/MM0_d N_XI9/NET18_XI9/XI142/MM0_g
+ N_XI9/XI142/NET043_XI9/XI142/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI140/MM0 N_WL<53>_XI9/XI140/MM0_d N_XI9/NET18_XI9/XI140/MM0_g
+ N_XI9/XI140/NET043_XI9/XI140/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI139/MM0 N_WL<52>_XI9/XI139/MM0_d N_XI9/NET18_XI9/XI139/MM0_g
+ N_XI9/XI139/NET043_XI9/XI139/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI144/MM0 N_WL<51>_XI9/XI144/MM0_d N_XI9/NET18_XI9/XI144/MM0_g
+ N_XI9/XI144/NET043_XI9/XI144/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI143/MM0 N_WL<50>_XI9/XI143/MM0_d N_XI9/NET18_XI9/XI143/MM0_g
+ N_XI9/XI143/NET043_XI9/XI143/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI145/MM0 N_WL<49>_XI9/XI145/MM0_d N_XI9/NET18_XI9/XI145/MM0_g
+ N_XI9/XI145/NET043_XI9/XI145/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI146/MM0 N_WL<48>_XI9/XI146/MM0_d N_XI9/NET18_XI9/XI146/MM0_g
+ N_XI9/XI146/NET043_XI9/XI146/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI125/MM0 N_WL<47>_XI9/XI125/MM0_d N_XI9/NET19_XI9/XI125/MM0_g
+ N_XI9/XI125/NET043_XI9/XI125/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI126/MM0 N_WL<46>_XI9/XI126/MM0_d N_XI9/NET19_XI9/XI126/MM0_g
+ N_XI9/XI126/NET043_XI9/XI126/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI124/MM0 N_WL<45>_XI9/XI124/MM0_d N_XI9/NET19_XI9/XI124/MM0_g
+ N_XI9/XI124/NET043_XI9/XI124/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI123/MM0 N_WL<44>_XI9/XI123/MM0_d N_XI9/NET19_XI9/XI123/MM0_g
+ N_XI9/XI123/NET043_XI9/XI123/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI128/MM0 N_WL<43>_XI9/XI128/MM0_d N_XI9/NET19_XI9/XI128/MM0_g
+ N_XI9/XI128/NET043_XI9/XI128/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI127/MM0 N_WL<42>_XI9/XI127/MM0_d N_XI9/NET19_XI9/XI127/MM0_g
+ N_XI9/XI127/NET043_XI9/XI127/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI129/MM0 N_WL<41>_XI9/XI129/MM0_d N_XI9/NET19_XI9/XI129/MM0_g
+ N_XI9/XI129/NET043_XI9/XI129/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI130/MM0 N_WL<40>_XI9/XI130/MM0_d N_XI9/NET19_XI9/XI130/MM0_g
+ N_XI9/XI130/NET043_XI9/XI130/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI120/MM0 N_WL<39>_XI9/XI120/MM0_d N_XI9/NET20_XI9/XI120/MM0_g
+ N_XI9/XI120/NET043_XI9/XI120/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI119/MM0 N_WL<38>_XI9/XI119/MM0_d N_XI9/NET20_XI9/XI119/MM0_g
+ N_XI9/XI119/NET043_XI9/XI119/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI121/MM0 N_WL<37>_XI9/XI121/MM0_d N_XI9/NET20_XI9/XI121/MM0_g
+ N_XI9/XI121/NET043_XI9/XI121/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI122/MM0 N_WL<36>_XI9/XI122/MM0_d N_XI9/NET20_XI9/XI122/MM0_g
+ N_XI9/XI122/NET043_XI9/XI122/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI117/MM0 N_WL<35>_XI9/XI117/MM0_d N_XI9/NET20_XI9/XI117/MM0_g
+ N_XI9/XI117/NET043_XI9/XI117/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI118/MM0 N_WL<34>_XI9/XI118/MM0_d N_XI9/NET20_XI9/XI118/MM0_g
+ N_XI9/XI118/NET043_XI9/XI118/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI116/MM0 N_WL<33>_XI9/XI116/MM0_d N_XI9/NET20_XI9/XI116/MM0_g
+ N_XI9/XI116/NET043_XI9/XI116/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI115/MM0 N_WL<32>_XI9/XI115/MM0_d N_XI9/NET20_XI9/XI115/MM0_g
+ N_XI9/XI115/NET043_XI9/XI115/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI104/MM0 N_WL<31>_XI9/XI104/MM0_d N_XI9/NET21_XI9/XI104/MM0_g
+ N_XI9/XI104/NET043_XI9/XI104/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI103/MM0 N_WL<30>_XI9/XI103/MM0_d N_XI9/NET21_XI9/XI103/MM0_g
+ N_XI9/XI103/NET043_XI9/XI103/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI105/MM0 N_WL<29>_XI9/XI105/MM0_d N_XI9/NET21_XI9/XI105/MM0_g
+ N_XI9/XI105/NET043_XI9/XI105/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI106/MM0 N_WL<28>_XI9/XI106/MM0_d N_XI9/NET21_XI9/XI106/MM0_g
+ N_XI9/XI106/NET043_XI9/XI106/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI101/MM0 N_WL<27>_XI9/XI101/MM0_d N_XI9/NET21_XI9/XI101/MM0_g
+ N_XI9/XI101/NET043_XI9/XI101/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI102/MM0 N_WL<26>_XI9/XI102/MM0_d N_XI9/NET21_XI9/XI102/MM0_g
+ N_XI9/XI102/NET043_XI9/XI102/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI100/MM0 N_WL<25>_XI9/XI100/MM0_d N_XI9/NET21_XI9/XI100/MM0_g
+ N_XI9/XI100/NET043_XI9/XI100/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI99/MM0 N_WL<24>_XI9/XI99/MM0_d N_XI9/NET21_XI9/XI99/MM0_g
+ N_XI9/XI99/NET043_XI9/XI99/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI109/MM0 N_WL<23>_XI9/XI109/MM0_d N_XI9/NET22_XI9/XI109/MM0_g
+ N_XI9/XI109/NET043_XI9/XI109/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI110/MM0 N_WL<22>_XI9/XI110/MM0_d N_XI9/NET22_XI9/XI110/MM0_g
+ N_XI9/XI110/NET043_XI9/XI110/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI108/MM0 N_WL<21>_XI9/XI108/MM0_d N_XI9/NET22_XI9/XI108/MM0_g
+ N_XI9/XI108/NET043_XI9/XI108/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI107/MM0 N_WL<20>_XI9/XI107/MM0_d N_XI9/NET22_XI9/XI107/MM0_g
+ N_XI9/XI107/NET043_XI9/XI107/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI112/MM0 N_WL<19>_XI9/XI112/MM0_d N_XI9/NET22_XI9/XI112/MM0_g
+ N_XI9/XI112/NET043_XI9/XI112/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI111/MM0 N_WL<18>_XI9/XI111/MM0_d N_XI9/NET22_XI9/XI111/MM0_g
+ N_XI9/XI111/NET043_XI9/XI111/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI113/MM0 N_WL<17>_XI9/XI113/MM0_d N_XI9/NET22_XI9/XI113/MM0_g
+ N_XI9/XI113/NET043_XI9/XI113/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI114/MM0 N_WL<16>_XI9/XI114/MM0_d N_XI9/NET22_XI9/XI114/MM0_g
+ N_XI9/XI114/NET043_XI9/XI114/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI93/MM0 N_WL<15>_XI9/XI93/MM0_d N_XI9/NET23_XI9/XI93/MM0_g
+ N_XI9/XI93/NET043_XI9/XI93/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI94/MM0 N_WL<14>_XI9/XI94/MM0_d N_XI9/NET23_XI9/XI94/MM0_g
+ N_XI9/XI94/NET043_XI9/XI94/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI92/MM0 N_WL<13>_XI9/XI92/MM0_d N_XI9/NET23_XI9/XI92/MM0_g
+ N_XI9/XI92/NET043_XI9/XI92/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI91/MM0 N_WL<12>_XI9/XI91/MM0_d N_XI9/NET23_XI9/XI91/MM0_g
+ N_XI9/XI91/NET043_XI9/XI91/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI96/MM0 N_WL<11>_XI9/XI96/MM0_d N_XI9/NET23_XI9/XI96/MM0_g
+ N_XI9/XI96/NET043_XI9/XI96/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI95/MM0 N_WL<10>_XI9/XI95/MM0_d N_XI9/NET23_XI9/XI95/MM0_g
+ N_XI9/XI95/NET043_XI9/XI95/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI97/MM0 N_WL<9>_XI9/XI97/MM0_d N_XI9/NET23_XI9/XI97/MM0_g
+ N_XI9/XI97/NET043_XI9/XI97/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI98/MM0 N_WL<8>_XI9/XI98/MM0_d N_XI9/NET23_XI9/XI98/MM0_g
+ N_XI9/XI98/NET043_XI9/XI98/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI88/MM0 N_WL<7>_XI9/XI88/MM0_d N_XI9/NET24_XI9/XI88/MM0_g
+ N_XI9/XI88/NET043_XI9/XI88/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI87/MM0 N_WL<6>_XI9/XI87/MM0_d N_XI9/NET24_XI9/XI87/MM0_g
+ N_XI9/XI87/NET043_XI9/XI87/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI89/MM0 N_WL<5>_XI9/XI89/MM0_d N_XI9/NET24_XI9/XI89/MM0_g
+ N_XI9/XI89/NET043_XI9/XI89/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI90/MM0 N_WL<4>_XI9/XI90/MM0_d N_XI9/NET24_XI9/XI90/MM0_g
+ N_XI9/XI90/NET043_XI9/XI90/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI85/MM0 N_WL<3>_XI9/XI85/MM0_d N_XI9/NET24_XI9/XI85/MM0_g
+ N_XI9/XI85/NET043_XI9/XI85/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI86/MM0 N_WL<2>_XI9/XI86/MM0_d N_XI9/NET24_XI9/XI86/MM0_g
+ N_XI9/XI86/NET043_XI9/XI86/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI84/MM0 N_WL<1>_XI9/XI84/MM0_d N_XI9/NET24_XI9/XI84/MM0_g
+ N_XI9/XI84/NET043_XI9/XI84/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI2/MM0 N_WL<0>_XI9/XI2/MM0_d N_XI9/NET24_XI9/XI2/MM0_g
+ N_XI9/XI2/NET043_XI9/XI2/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI136/MM10 N_XI9/XI136/NET043_XI9/XI136/MM10_d N_XI9/NET4_XI9/XI136/MM10_g
+ N_VDD_XI9/XI136/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI135/MM10 N_XI9/XI135/NET043_XI9/XI135/MM10_d N_XI9/NET5_XI9/XI135/MM10_g
+ N_VDD_XI9/XI135/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI137/MM10 N_XI9/XI137/NET043_XI9/XI137/MM10_d N_XI9/NET6_XI9/XI137/MM10_g
+ N_VDD_XI9/XI137/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI138/MM10 N_XI9/XI138/NET043_XI9/XI138/MM10_d N_XI9/NET7_XI9/XI138/MM10_g
+ N_VDD_XI9/XI138/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI133/MM10 N_XI9/XI133/NET043_XI9/XI133/MM10_d N_XI9/NET8_XI9/XI133/MM10_g
+ N_VDD_XI9/XI133/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI134/MM10 N_XI9/XI134/NET043_XI9/XI134/MM10_d N_XI9/NET9_XI9/XI134/MM10_g
+ N_VDD_XI9/XI134/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI132/MM10 N_XI9/XI132/NET043_XI9/XI132/MM10_d N_XI9/NET10_XI9/XI132/MM10_g
+ N_VDD_XI9/XI132/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI131/MM10 N_XI9/XI131/NET043_XI9/XI131/MM10_d N_XI9/NET11_XI9/XI131/MM10_g
+ N_VDD_XI9/XI131/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI141/MM10 N_XI9/XI141/NET043_XI9/XI141/MM10_d N_XI9/NET4_XI9/XI141/MM10_g
+ N_VDD_XI9/XI141/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI142/MM10 N_XI9/XI142/NET043_XI9/XI142/MM10_d N_XI9/NET5_XI9/XI142/MM10_g
+ N_VDD_XI9/XI142/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI140/MM10 N_XI9/XI140/NET043_XI9/XI140/MM10_d N_XI9/NET6_XI9/XI140/MM10_g
+ N_VDD_XI9/XI140/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI139/MM10 N_XI9/XI139/NET043_XI9/XI139/MM10_d N_XI9/NET7_XI9/XI139/MM10_g
+ N_VDD_XI9/XI139/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI144/MM10 N_XI9/XI144/NET043_XI9/XI144/MM10_d N_XI9/NET8_XI9/XI144/MM10_g
+ N_VDD_XI9/XI144/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI143/MM10 N_XI9/XI143/NET043_XI9/XI143/MM10_d N_XI9/NET9_XI9/XI143/MM10_g
+ N_VDD_XI9/XI143/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI145/MM10 N_XI9/XI145/NET043_XI9/XI145/MM10_d N_XI9/NET10_XI9/XI145/MM10_g
+ N_VDD_XI9/XI145/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI146/MM10 N_XI9/XI146/NET043_XI9/XI146/MM10_d N_XI9/NET11_XI9/XI146/MM10_g
+ N_VDD_XI9/XI146/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI125/MM10 N_XI9/XI125/NET043_XI9/XI125/MM10_d N_XI9/NET4_XI9/XI125/MM10_g
+ N_VDD_XI9/XI125/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI126/MM10 N_XI9/XI126/NET043_XI9/XI126/MM10_d N_XI9/NET5_XI9/XI126/MM10_g
+ N_VDD_XI9/XI126/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI124/MM10 N_XI9/XI124/NET043_XI9/XI124/MM10_d N_XI9/NET6_XI9/XI124/MM10_g
+ N_VDD_XI9/XI124/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI123/MM10 N_XI9/XI123/NET043_XI9/XI123/MM10_d N_XI9/NET7_XI9/XI123/MM10_g
+ N_VDD_XI9/XI123/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI128/MM10 N_XI9/XI128/NET043_XI9/XI128/MM10_d N_XI9/NET8_XI9/XI128/MM10_g
+ N_VDD_XI9/XI128/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI127/MM10 N_XI9/XI127/NET043_XI9/XI127/MM10_d N_XI9/NET9_XI9/XI127/MM10_g
+ N_VDD_XI9/XI127/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI129/MM10 N_XI9/XI129/NET043_XI9/XI129/MM10_d N_XI9/NET10_XI9/XI129/MM10_g
+ N_VDD_XI9/XI129/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI130/MM10 N_XI9/XI130/NET043_XI9/XI130/MM10_d N_XI9/NET11_XI9/XI130/MM10_g
+ N_VDD_XI9/XI130/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI120/MM10 N_XI9/XI120/NET043_XI9/XI120/MM10_d N_XI9/NET4_XI9/XI120/MM10_g
+ N_VDD_XI9/XI120/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI119/MM10 N_XI9/XI119/NET043_XI9/XI119/MM10_d N_XI9/NET5_XI9/XI119/MM10_g
+ N_VDD_XI9/XI119/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI121/MM10 N_XI9/XI121/NET043_XI9/XI121/MM10_d N_XI9/NET6_XI9/XI121/MM10_g
+ N_VDD_XI9/XI121/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI122/MM10 N_XI9/XI122/NET043_XI9/XI122/MM10_d N_XI9/NET7_XI9/XI122/MM10_g
+ N_VDD_XI9/XI122/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI117/MM10 N_XI9/XI117/NET043_XI9/XI117/MM10_d N_XI9/NET8_XI9/XI117/MM10_g
+ N_VDD_XI9/XI117/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI118/MM10 N_XI9/XI118/NET043_XI9/XI118/MM10_d N_XI9/NET9_XI9/XI118/MM10_g
+ N_VDD_XI9/XI118/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI116/MM10 N_XI9/XI116/NET043_XI9/XI116/MM10_d N_XI9/NET10_XI9/XI116/MM10_g
+ N_VDD_XI9/XI116/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI115/MM10 N_XI9/XI115/NET043_XI9/XI115/MM10_d N_XI9/NET11_XI9/XI115/MM10_g
+ N_VDD_XI9/XI115/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI104/MM10 N_XI9/XI104/NET043_XI9/XI104/MM10_d N_XI9/NET4_XI9/XI104/MM10_g
+ N_VDD_XI9/XI104/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI103/MM10 N_XI9/XI103/NET043_XI9/XI103/MM10_d N_XI9/NET5_XI9/XI103/MM10_g
+ N_VDD_XI9/XI103/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI105/MM10 N_XI9/XI105/NET043_XI9/XI105/MM10_d N_XI9/NET6_XI9/XI105/MM10_g
+ N_VDD_XI9/XI105/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI106/MM10 N_XI9/XI106/NET043_XI9/XI106/MM10_d N_XI9/NET7_XI9/XI106/MM10_g
+ N_VDD_XI9/XI106/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI101/MM10 N_XI9/XI101/NET043_XI9/XI101/MM10_d N_XI9/NET8_XI9/XI101/MM10_g
+ N_VDD_XI9/XI101/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI102/MM10 N_XI9/XI102/NET043_XI9/XI102/MM10_d N_XI9/NET9_XI9/XI102/MM10_g
+ N_VDD_XI9/XI102/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI100/MM10 N_XI9/XI100/NET043_XI9/XI100/MM10_d N_XI9/NET10_XI9/XI100/MM10_g
+ N_VDD_XI9/XI100/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI99/MM10 N_XI9/XI99/NET043_XI9/XI99/MM10_d N_XI9/NET11_XI9/XI99/MM10_g
+ N_VDD_XI9/XI99/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI109/MM10 N_XI9/XI109/NET043_XI9/XI109/MM10_d N_XI9/NET4_XI9/XI109/MM10_g
+ N_VDD_XI9/XI109/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI110/MM10 N_XI9/XI110/NET043_XI9/XI110/MM10_d N_XI9/NET5_XI9/XI110/MM10_g
+ N_VDD_XI9/XI110/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI108/MM10 N_XI9/XI108/NET043_XI9/XI108/MM10_d N_XI9/NET6_XI9/XI108/MM10_g
+ N_VDD_XI9/XI108/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI107/MM10 N_XI9/XI107/NET043_XI9/XI107/MM10_d N_XI9/NET7_XI9/XI107/MM10_g
+ N_VDD_XI9/XI107/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI112/MM10 N_XI9/XI112/NET043_XI9/XI112/MM10_d N_XI9/NET8_XI9/XI112/MM10_g
+ N_VDD_XI9/XI112/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI111/MM10 N_XI9/XI111/NET043_XI9/XI111/MM10_d N_XI9/NET9_XI9/XI111/MM10_g
+ N_VDD_XI9/XI111/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI113/MM10 N_XI9/XI113/NET043_XI9/XI113/MM10_d N_XI9/NET10_XI9/XI113/MM10_g
+ N_VDD_XI9/XI113/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI114/MM10 N_XI9/XI114/NET043_XI9/XI114/MM10_d N_XI9/NET11_XI9/XI114/MM10_g
+ N_VDD_XI9/XI114/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI93/MM10 N_XI9/XI93/NET043_XI9/XI93/MM10_d N_XI9/NET4_XI9/XI93/MM10_g
+ N_VDD_XI9/XI93/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI94/MM10 N_XI9/XI94/NET043_XI9/XI94/MM10_d N_XI9/NET5_XI9/XI94/MM10_g
+ N_VDD_XI9/XI94/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI92/MM10 N_XI9/XI92/NET043_XI9/XI92/MM10_d N_XI9/NET6_XI9/XI92/MM10_g
+ N_VDD_XI9/XI92/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI91/MM10 N_XI9/XI91/NET043_XI9/XI91/MM10_d N_XI9/NET7_XI9/XI91/MM10_g
+ N_VDD_XI9/XI91/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI96/MM10 N_XI9/XI96/NET043_XI9/XI96/MM10_d N_XI9/NET8_XI9/XI96/MM10_g
+ N_VDD_XI9/XI96/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI95/MM10 N_XI9/XI95/NET043_XI9/XI95/MM10_d N_XI9/NET9_XI9/XI95/MM10_g
+ N_VDD_XI9/XI95/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI97/MM10 N_XI9/XI97/NET043_XI9/XI97/MM10_d N_XI9/NET10_XI9/XI97/MM10_g
+ N_VDD_XI9/XI97/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI98/MM10 N_XI9/XI98/NET043_XI9/XI98/MM10_d N_XI9/NET11_XI9/XI98/MM10_g
+ N_VDD_XI9/XI98/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI88/MM10 N_XI9/XI88/NET043_XI9/XI88/MM10_d N_XI9/NET4_XI9/XI88/MM10_g
+ N_VDD_XI9/XI88/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI87/MM10 N_XI9/XI87/NET043_XI9/XI87/MM10_d N_XI9/NET5_XI9/XI87/MM10_g
+ N_VDD_XI9/XI87/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI89/MM10 N_XI9/XI89/NET043_XI9/XI89/MM10_d N_XI9/NET6_XI9/XI89/MM10_g
+ N_VDD_XI9/XI89/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI90/MM10 N_XI9/XI90/NET043_XI9/XI90/MM10_d N_XI9/NET7_XI9/XI90/MM10_g
+ N_VDD_XI9/XI90/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI85/MM10 N_XI9/XI85/NET043_XI9/XI85/MM10_d N_XI9/NET8_XI9/XI85/MM10_g
+ N_VDD_XI9/XI85/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI86/MM10 N_XI9/XI86/NET043_XI9/XI86/MM10_d N_XI9/NET9_XI9/XI86/MM10_g
+ N_VDD_XI9/XI86/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI84/MM10 N_XI9/XI84/NET043_XI9/XI84/MM10_d N_XI9/NET10_XI9/XI84/MM10_g
+ N_VDD_XI9/XI84/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9/XI2/MM10 N_XI9/XI2/NET043_XI9/XI2/MM10_d N_XI9/NET11_XI9/XI2/MM10_g
+ N_VDD_XI9/XI2/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI13/MM8 N_BL<0>_XI13/MM8_d N_CLK_XI13/MM8_g N_VDD_XI13/MM8_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI16/XI21/XI1/MM6 N_XI16/XI21/NET40_XI16/XI21/XI1/MM6_d
+ N_YOUT<1>_XI16/XI21/XI1/MM6_g N_VDD_XI16/XI21/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI16/XI21/MM0 N_BL<1>_XI16/XI21/MM0_d N_YOUT<1>_XI16/XI21/MM0_g
+ N_DL<0>_XI16/XI21/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI22/XI1/MM6 N_XI16/XI22/NET40_XI16/XI22/XI1/MM6_d
+ N_YOUT<0>_XI16/XI22/XI1/MM6_g N_VDD_XI16/XI22/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI22/MM0 N_BL<0>_XI16/XI22/MM0_d N_YOUT<0>_XI16/XI22/MM0_g
+ N_DL<0>_XI16/XI22/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM9 N_BL<1>_XI13/MM9_d N_CLK_XI13/MM9_g N_VDD_XI13/MM9_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI13/MM10 N_BL<2>_XI13/MM10_d N_CLK_XI13/MM10_g N_VDD_XI13/MM10_s
+ N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXI16/XI19/XI1/MM6 N_XI16/XI19/NET40_XI16/XI19/XI1/MM6_d
+ N_YOUT<3>_XI16/XI19/XI1/MM6_g N_VDD_XI16/XI19/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI16/XI19/MM0 N_BL<3>_XI16/XI19/MM0_d N_YOUT<3>_XI16/XI19/MM0_g
+ N_DL<0>_XI16/XI19/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI20/XI1/MM6 N_XI16/XI20/NET40_XI16/XI20/XI1/MM6_d
+ N_YOUT<2>_XI16/XI20/XI1/MM6_g N_VDD_XI16/XI20/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI20/MM0 N_BL<2>_XI16/XI20/MM0_d N_YOUT<2>_XI16/XI20/MM0_g
+ N_DL<0>_XI16/XI20/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM11 N_BL<3>_XI13/MM11_d N_CLK_XI13/MM11_g N_VDD_XI13/MM11_s
+ N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXI13/MM12 N_BL<4>_XI13/MM12_d N_CLK_XI13/MM12_g N_VDD_XI13/MM12_s
+ N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXI16/XI16/XI1/MM6 N_XI16/XI16/NET40_XI16/XI16/XI1/MM6_d
+ N_YOUT<5>_XI16/XI16/XI1/MM6_g N_VDD_XI16/XI16/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI16/XI16/MM0 N_BL<5>_XI16/XI16/MM0_d N_YOUT<5>_XI16/XI16/MM0_g
+ N_DL<0>_XI16/XI16/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI15/XI1/MM6 N_XI16/XI15/NET40_XI16/XI15/XI1/MM6_d
+ N_YOUT<4>_XI16/XI15/XI1/MM6_g N_VDD_XI16/XI15/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI15/MM0 N_BL<4>_XI16/XI15/MM0_d N_YOUT<4>_XI16/XI15/MM0_g
+ N_DL<0>_XI16/XI15/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM13 N_BL<5>_XI13/MM13_d N_CLK_XI13/MM13_g N_VDD_XI13/MM13_s
+ N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXI13/MM14 N_BL<6>_XI13/MM14_d N_CLK_XI13/MM14_g N_VDD_XI13/MM14_s
+ N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXI16/XI18/XI1/MM6 N_XI16/XI18/NET40_XI16/XI18/XI1/MM6_d
+ N_YOUT<7>_XI16/XI18/XI1/MM6_g N_VDD_XI16/XI18/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI16/XI18/MM0 N_BL<7>_XI16/XI18/MM0_d N_YOUT<7>_XI16/XI18/MM0_g
+ N_DL<0>_XI16/XI18/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI17/XI1/MM6 N_XI16/XI17/NET40_XI16/XI17/XI1/MM6_d
+ N_YOUT<6>_XI16/XI17/XI1/MM6_g N_VDD_XI16/XI17/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI16/XI17/MM0 N_BL<6>_XI16/XI17/MM0_d N_YOUT<6>_XI16/XI17/MM0_g
+ N_DL<0>_XI16/XI17/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM15 N_BL<7>_XI13/MM15_d N_CLK_XI13/MM15_g N_VDD_XI13/MM15_s
+ N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXI13/MM7 N_BL<8>_XI13/MM7_d N_CLK_XI13/MM7_g N_VDD_XI13/MM7_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI17/XI21/XI1/MM6 N_XI17/XI21/NET40_XI17/XI21/XI1/MM6_d
+ N_YOUT<1>_XI17/XI21/XI1/MM6_g N_VDD_XI17/XI21/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI17/XI21/MM0 N_BL<9>_XI17/XI21/MM0_d N_YOUT<1>_XI17/XI21/MM0_g
+ N_DL<1>_XI17/XI21/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI22/XI1/MM6 N_XI17/XI22/NET40_XI17/XI22/XI1/MM6_d
+ N_YOUT<0>_XI17/XI22/XI1/MM6_g N_VDD_XI17/XI22/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI22/MM0 N_BL<8>_XI17/XI22/MM0_d N_YOUT<0>_XI17/XI22/MM0_g
+ N_DL<1>_XI17/XI22/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM6 N_BL<9>_XI13/MM6_d N_CLK_XI13/MM6_g N_VDD_XI13/MM6_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI13/MM5 N_BL<10>_XI13/MM5_d N_CLK_XI13/MM5_g N_VDD_XI13/MM5_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI17/XI19/XI1/MM6 N_XI17/XI19/NET40_XI17/XI19/XI1/MM6_d
+ N_YOUT<3>_XI17/XI19/XI1/MM6_g N_VDD_XI17/XI19/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI17/XI19/MM0 N_BL<11>_XI17/XI19/MM0_d N_YOUT<3>_XI17/XI19/MM0_g
+ N_DL<1>_XI17/XI19/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI20/XI1/MM6 N_XI17/XI20/NET40_XI17/XI20/XI1/MM6_d
+ N_YOUT<2>_XI17/XI20/XI1/MM6_g N_VDD_XI17/XI20/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI20/MM0 N_BL<10>_XI17/XI20/MM0_d N_YOUT<2>_XI17/XI20/MM0_g
+ N_DL<1>_XI17/XI20/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM4 N_BL<11>_XI13/MM4_d N_CLK_XI13/MM4_g N_VDD_XI13/MM4_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI13/MM3 N_BL<12>_XI13/MM3_d N_CLK_XI13/MM3_g N_VDD_XI13/MM3_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI17/XI16/XI1/MM6 N_XI17/XI16/NET40_XI17/XI16/XI1/MM6_d
+ N_YOUT<5>_XI17/XI16/XI1/MM6_g N_VDD_XI17/XI16/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI17/XI16/MM0 N_BL<13>_XI17/XI16/MM0_d N_YOUT<5>_XI17/XI16/MM0_g
+ N_DL<1>_XI17/XI16/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI15/XI1/MM6 N_XI17/XI15/NET40_XI17/XI15/XI1/MM6_d
+ N_YOUT<4>_XI17/XI15/XI1/MM6_g N_VDD_XI17/XI15/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI15/MM0 N_BL<12>_XI17/XI15/MM0_d N_YOUT<4>_XI17/XI15/MM0_g
+ N_DL<1>_XI17/XI15/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM2 N_BL<13>_XI13/MM2_d N_CLK_XI13/MM2_g N_VDD_XI13/MM2_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI13/MM1 N_BL<14>_XI13/MM1_d N_CLK_XI13/MM1_g N_VDD_XI13/MM1_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI17/XI18/XI1/MM6 N_XI17/XI18/NET40_XI17/XI18/XI1/MM6_d
+ N_YOUT<7>_XI17/XI18/XI1/MM6_g N_VDD_XI17/XI18/XI1/MM6_s
+ N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI17/XI18/MM0 N_BL<15>_XI17/XI18/MM0_d N_YOUT<7>_XI17/XI18/MM0_g
+ N_DL<1>_XI17/XI18/MM0_s N_VDD_XI16/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI17/XI1/MM6 N_XI17/XI17/NET40_XI17/XI17/XI1/MM6_d
+ N_YOUT<6>_XI17/XI17/XI1/MM6_g N_VDD_XI17/XI17/XI1/MM6_s N_VDD_XI13/MM8_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI17/XI17/MM0 N_BL<14>_XI17/XI17/MM0_d N_YOUT<6>_XI17/XI17/MM0_g
+ N_DL<1>_XI17/XI17/MM0_s N_VDD_XI13/MM8_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI13/MM0 N_BL<15>_XI13/MM0_d N_CLK_XI13/MM0_g N_VDD_XI13/MM0_s N_VDD_XI13/MM8_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07
mXI27/MM16 N_XI27/NET093_XI27/MM16_d N_DL<0>_XI27/MM16_g
+ N_XI27/NET096_XI27/MM16_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI27/MM19 N_XI27/NET096_XI27/MM19_d N_SAEN_XI27/MM19_g N_VSS_XI27/MM19_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06
+ PS=5.1e-07
mXI27/MM15 N_SO<0>_XI27/MM15_d N_DOUT<0>_XI27/MM15_g N_XI27/NET093_XI27/MM15_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI27/MM19@4 N_XI27/NET096_XI27/MM19@4_d N_SAEN_XI27/MM19@4_g
+ N_VSS_XI27/MM19@4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXI27/MM19@3 N_XI27/NET096_XI27/MM19@3_d N_SAEN_XI27/MM19@3_g
+ N_VSS_XI27/MM19@3_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXI27/MM17 N_DOUT<0>_XI27/MM17_d N_SO<0>_XI27/MM17_g N_XI27/NET089_XI27/MM17_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI27/MM19@2 N_XI27/NET096_XI27/MM19@2_d N_SAEN_XI27/MM19@2_g
+ N_VSS_XI27/MM19@2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXI27/MM18 N_XI27/NET089_XI27/MM18_d N_VREF_XI27/MM18_g
+ N_XI27/NET096_XI27/MM18_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI27/MM11 N_SO<0>_XI27/MM11_d N_SAEN_XI27/MM11_g N_VDD_XI27/MM11_s
+ N_VDD_XI27/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI27/MM12 N_SO<0>_XI27/MM12_d N_DOUT<0>_XI27/MM12_g N_VDD_XI27/MM12_s
+ N_VDD_XI27/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI27/MM13 N_DOUT<0>_XI27/MM13_d N_SO<0>_XI27/MM13_g N_VDD_XI27/MM13_s
+ N_VDD_XI27/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI27/MM9 N_DOUT<0>_XI27/MM9_d N_SAEN_XI27/MM9_g N_VDD_XI27/MM9_s
+ N_VDD_XI27/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI28/MM16 N_XI28/NET093_XI28/MM16_d N_DL<1>_XI28/MM16_g
+ N_XI28/NET096_XI28/MM16_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI28/MM19 N_XI28/NET096_XI28/MM19_d N_SAEN_XI28/MM19_g N_VSS_XI28/MM19_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06
+ PS=5.1e-07
mXI28/MM15 N_SO<1>_XI28/MM15_d N_DOUT<1>_XI28/MM15_g N_XI28/NET093_XI28/MM15_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI28/MM19@4 N_XI28/NET096_XI28/MM19@4_d N_SAEN_XI28/MM19@4_g
+ N_VSS_XI28/MM19@4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXI28/MM19@3 N_XI28/NET096_XI28/MM19@3_d N_SAEN_XI28/MM19@3_g
+ N_VSS_XI28/MM19@3_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXI28/MM17 N_DOUT<1>_XI28/MM17_d N_SO<1>_XI28/MM17_g N_XI28/NET089_XI28/MM17_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI28/MM19@2 N_XI28/NET096_XI28/MM19@2_d N_SAEN_XI28/MM19@2_g
+ N_VSS_XI28/MM19@2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXI28/MM18 N_XI28/NET089_XI28/MM18_d N_VREF_XI28/MM18_g
+ N_XI28/NET096_XI28/MM18_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI28/MM11 N_SO<1>_XI28/MM11_d N_SAEN_XI28/MM11_g N_VDD_XI28/MM11_s
+ N_VDD_XI28/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI28/MM12 N_SO<1>_XI28/MM12_d N_DOUT<1>_XI28/MM12_g N_VDD_XI28/MM12_s
+ N_VDD_XI28/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI28/MM13 N_DOUT<1>_XI28/MM13_d N_SO<1>_XI28/MM13_g N_VDD_XI28/MM13_s
+ N_VDD_XI28/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI28/MM9 N_DOUT<1>_XI28/MM9_d N_SAEN_XI28/MM9_g N_VDD_XI28/MM9_s
+ N_VDD_XI28/MM11_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI29/XI44/MM10 N_XI29/NET0145_XI29/XI44/MM10_d N_CLK_XI29/XI44/MM10_g
+ N_VSS_XI29/XI44/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI44/MM6 N_XI29/NET0145_XI29/XI44/MM6_d N_CLK_XI29/XI44/MM6_g
+ N_VDD_XI29/XI44/MM6_s N_VDD_XI29/XI44/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI50/XI5/MM10 N_XI29/XI50/NET14_XI29/XI50/XI5/MM10_d
+ N_XI29/NET0146_XI29/XI50/XI5/MM10_g N_VSS_XI29/XI50/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI50/XI5/MM6 N_XI29/XI50/NET14_XI29/XI50/XI5/MM6_d
+ N_XI29/NET0146_XI29/XI50/XI5/MM6_g N_VDD_XI29/XI50/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI42/MM5 N_XI29/XI42/NET44_XI29/XI42/MM5_d N_XI29/NET101_XI29/XI42/MM5_g
+ N_VSS_XI29/XI42/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI29/XI42/MM4 N_XI29/XI42/NET067_XI29/XI42/MM4_d N_CLK_XI29/XI42/MM4_g
+ N_XI29/XI42/NET44_XI29/XI42/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI29/XI42/MM0 N_XI29/XI42/NET067_XI29/XI42/MM0_d N_XI29/NET101_XI29/XI42/MM0_g
+ N_VDD_XI29/XI42/MM0_s N_VDD_XI29/XI42/MM9_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI29/XI42/MM1 N_XI29/XI42/NET067_XI29/XI42/MM1_d N_CLK_XI29/XI42/MM1_g
+ N_VDD_XI29/XI42/MM1_s N_VDD_XI29/XI42/MM9_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI29/XI42/MM10 N_WLEN_XI29/XI42/MM10_d N_XI29/XI42/NET067_XI29/XI42/MM10_g
+ N_VSS_XI29/XI42/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI42/MM9 N_WLEN_XI29/XI42/MM9_d N_XI29/XI42/NET067_XI29/XI42/MM9_g
+ N_VDD_XI29/XI42/MM9_s N_VDD_XI29/XI42/MM9_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI43/MM5 N_XI29/XI43/NET44_XI29/XI43/MM5_d N_XI29/NET0134_XI29/XI43/MM5_g
+ N_VSS_XI29/XI43/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI29/XI43/MM4 N_XI29/XI43/NET067_XI29/XI43/MM4_d N_CLK_XI29/XI43/MM4_g
+ N_XI29/XI43/NET44_XI29/XI43/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI29/XI43/MM0 N_XI29/XI43/NET067_XI29/XI43/MM0_d N_XI29/NET0134_XI29/XI43/MM0_g
+ N_VDD_XI29/XI43/MM0_s N_VDD_XI29/XI43/MM9_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI29/XI43/MM1 N_XI29/XI43/NET067_XI29/XI43/MM1_d N_CLK_XI29/XI43/MM1_g
+ N_VDD_XI29/XI43/MM1_s N_VDD_XI29/XI43/MM9_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI29/XI43/MM10 N_SAEN_XI29/XI43/MM10_d N_XI29/XI43/NET067_XI29/XI43/MM10_g
+ N_VSS_XI29/XI43/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI43/MM9 N_SAEN_XI29/XI43/MM9_d N_XI29/XI43/NET067_XI29/XI43/MM9_g
+ N_VDD_XI29/XI43/MM9_s N_VDD_XI29/XI43/MM9_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI26/XI3/MM11 N_XI26/XI3/NET030_XI26/XI3/MM11_d N_VDD_XI26/XI3/MM11_g
+ N_VSS_XI26/XI3/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI3/MM6 N_XI26/XI3/NET40_XI26/XI3/MM6_d N_Y_SEL<2>_XI26/XI3/MM6_g
+ N_XI26/XI3/NET030_XI26/XI3/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI3/MM5 N_XI26/XI3/NET44_XI26/XI3/MM5_d N_Y_SEL<1>_XI26/XI3/MM5_g
+ N_XI26/XI3/NET40_XI26/XI3/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI3/MM4 N_YOUT<3>_XI26/XI3/MM4_d N_XI26/NET0158_XI26/XI3/MM4_g
+ N_XI26/XI3/NET44_XI26/XI3/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI2/MM11 N_XI26/XI2/NET030_XI26/XI2/MM11_d N_VDD_XI26/XI2/MM11_g
+ N_VSS_XI26/XI2/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI2/MM6 N_XI26/XI2/NET40_XI26/XI2/MM6_d N_XI26/NET0116_XI26/XI2/MM6_g
+ N_XI26/XI2/NET030_XI26/XI2/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI2/MM5 N_XI26/XI2/NET44_XI26/XI2/MM5_d N_Y_SEL<1>_XI26/XI2/MM5_g
+ N_XI26/XI2/NET40_XI26/XI2/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI2/MM4 N_YOUT<2>_XI26/XI2/MM4_d N_XI26/NET0158_XI26/XI2/MM4_g
+ N_XI26/XI2/NET44_XI26/XI2/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI1/MM11 N_XI26/XI1/NET030_XI26/XI1/MM11_d N_VDD_XI26/XI1/MM11_g
+ N_VSS_XI26/XI1/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI1/MM6 N_XI26/XI1/NET40_XI26/XI1/MM6_d N_Y_SEL<2>_XI26/XI1/MM6_g
+ N_XI26/XI1/NET030_XI26/XI1/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI1/MM5 N_XI26/XI1/NET44_XI26/XI1/MM5_d N_XI26/NET0105_XI26/XI1/MM5_g
+ N_XI26/XI1/NET40_XI26/XI1/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI1/MM4 N_YOUT<1>_XI26/XI1/MM4_d N_XI26/NET0158_XI26/XI1/MM4_g
+ N_XI26/XI1/NET44_XI26/XI1/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI0/MM11 N_XI26/XI0/NET030_XI26/XI0/MM11_d N_VDD_XI26/XI0/MM11_g
+ N_VSS_XI26/XI0/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI0/MM6 N_XI26/XI0/NET40_XI26/XI0/MM6_d N_XI26/NET0116_XI26/XI0/MM6_g
+ N_XI26/XI0/NET030_XI26/XI0/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI0/MM5 N_XI26/XI0/NET44_XI26/XI0/MM5_d N_XI26/NET0105_XI26/XI0/MM5_g
+ N_XI26/XI0/NET40_XI26/XI0/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI0/MM4 N_YOUT<0>_XI26/XI0/MM4_d N_XI26/NET0158_XI26/XI0/MM4_g
+ N_XI26/XI0/NET44_XI26/XI0/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI7/MM11 N_XI26/XI7/NET030_XI26/XI7/MM11_d N_VDD_XI26/XI7/MM11_g
+ N_VSS_XI26/XI7/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI7/MM6 N_XI26/XI7/NET40_XI26/XI7/MM6_d N_Y_SEL<2>_XI26/XI7/MM6_g
+ N_XI26/XI7/NET030_XI26/XI7/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI7/MM5 N_XI26/XI7/NET44_XI26/XI7/MM5_d N_Y_SEL<1>_XI26/XI7/MM5_g
+ N_XI26/XI7/NET40_XI26/XI7/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI7/MM4 N_YOUT<7>_XI26/XI7/MM4_d N_Y_SEL<0>_XI26/XI7/MM4_g
+ N_XI26/XI7/NET44_XI26/XI7/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI6/MM11 N_XI26/XI6/NET030_XI26/XI6/MM11_d N_VDD_XI26/XI6/MM11_g
+ N_VSS_XI26/XI6/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI6/MM6 N_XI26/XI6/NET40_XI26/XI6/MM6_d N_XI26/NET0116_XI26/XI6/MM6_g
+ N_XI26/XI6/NET030_XI26/XI6/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI6/MM5 N_XI26/XI6/NET44_XI26/XI6/MM5_d N_Y_SEL<1>_XI26/XI6/MM5_g
+ N_XI26/XI6/NET40_XI26/XI6/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI6/MM4 N_YOUT<6>_XI26/XI6/MM4_d N_Y_SEL<0>_XI26/XI6/MM4_g
+ N_XI26/XI6/NET44_XI26/XI6/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI5/MM11 N_XI26/XI5/NET030_XI26/XI5/MM11_d N_VDD_XI26/XI5/MM11_g
+ N_VSS_XI26/XI5/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI5/MM6 N_XI26/XI5/NET40_XI26/XI5/MM6_d N_Y_SEL<2>_XI26/XI5/MM6_g
+ N_XI26/XI5/NET030_XI26/XI5/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI5/MM5 N_XI26/XI5/NET44_XI26/XI5/MM5_d N_XI26/NET0105_XI26/XI5/MM5_g
+ N_XI26/XI5/NET40_XI26/XI5/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI5/MM4 N_YOUT<5>_XI26/XI5/MM4_d N_Y_SEL<0>_XI26/XI5/MM4_g
+ N_XI26/XI5/NET44_XI26/XI5/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI4/MM11 N_XI26/XI4/NET030_XI26/XI4/MM11_d N_VDD_XI26/XI4/MM11_g
+ N_VSS_XI26/XI4/MM11_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI4/MM6 N_XI26/XI4/NET40_XI26/XI4/MM6_d N_XI26/NET0116_XI26/XI4/MM6_g
+ N_XI26/XI4/NET030_XI26/XI4/MM6_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI4/MM5 N_XI26/XI4/NET44_XI26/XI4/MM5_d N_XI26/NET0105_XI26/XI4/MM5_g
+ N_XI26/XI4/NET40_XI26/XI4/MM5_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI4/MM4 N_YOUT<4>_XI26/XI4/MM4_d N_Y_SEL<0>_XI26/XI4/MM4_g
+ N_XI26/XI4/NET44_XI26/XI4/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI26/XI3/MM12 N_YOUT<3>_XI26/XI3/MM12_d N_VDD_XI26/XI3/MM12_g
+ N_VDD_XI26/XI3/MM12_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI3/MM2 N_YOUT<3>_XI26/XI3/MM2_d N_Y_SEL<2>_XI26/XI3/MM2_g
+ N_VDD_XI26/XI3/MM2_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI3/MM0 N_YOUT<3>_XI26/XI3/MM0_d N_Y_SEL<1>_XI26/XI3/MM0_g
+ N_VDD_XI26/XI3/MM0_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI3/MM10 N_YOUT<3>_XI26/XI3/MM10_d N_XI26/NET0158_XI26/XI3/MM10_g
+ N_VDD_XI26/XI3/MM10_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI2/MM12 N_YOUT<2>_XI26/XI2/MM12_d N_VDD_XI26/XI2/MM12_g
+ N_VDD_XI26/XI2/MM12_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI2/MM2 N_YOUT<2>_XI26/XI2/MM2_d N_XI26/NET0116_XI26/XI2/MM2_g
+ N_VDD_XI26/XI2/MM2_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI2/MM0 N_YOUT<2>_XI26/XI2/MM0_d N_Y_SEL<1>_XI26/XI2/MM0_g
+ N_VDD_XI26/XI2/MM0_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI2/MM10 N_YOUT<2>_XI26/XI2/MM10_d N_XI26/NET0158_XI26/XI2/MM10_g
+ N_VDD_XI26/XI2/MM10_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI1/MM12 N_YOUT<1>_XI26/XI1/MM12_d N_VDD_XI26/XI1/MM12_g
+ N_VDD_XI26/XI1/MM12_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI1/MM2 N_YOUT<1>_XI26/XI1/MM2_d N_Y_SEL<2>_XI26/XI1/MM2_g
+ N_VDD_XI26/XI1/MM2_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI1/MM0 N_YOUT<1>_XI26/XI1/MM0_d N_XI26/NET0105_XI26/XI1/MM0_g
+ N_VDD_XI26/XI1/MM0_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI1/MM10 N_YOUT<1>_XI26/XI1/MM10_d N_XI26/NET0158_XI26/XI1/MM10_g
+ N_VDD_XI26/XI1/MM10_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI0/MM12 N_YOUT<0>_XI26/XI0/MM12_d N_VDD_XI26/XI0/MM12_g
+ N_VDD_XI26/XI0/MM12_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI0/MM2 N_YOUT<0>_XI26/XI0/MM2_d N_XI26/NET0116_XI26/XI0/MM2_g
+ N_VDD_XI26/XI0/MM2_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI0/MM0 N_YOUT<0>_XI26/XI0/MM0_d N_XI26/NET0105_XI26/XI0/MM0_g
+ N_VDD_XI26/XI0/MM0_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI0/MM10 N_YOUT<0>_XI26/XI0/MM10_d N_XI26/NET0158_XI26/XI0/MM10_g
+ N_VDD_XI26/XI0/MM10_s N_VDD_XI26/XI3/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI7/MM12 N_YOUT<7>_XI26/XI7/MM12_d N_VDD_XI26/XI7/MM12_g
+ N_VDD_XI26/XI7/MM12_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI7/MM2 N_YOUT<7>_XI26/XI7/MM2_d N_Y_SEL<2>_XI26/XI7/MM2_g
+ N_VDD_XI26/XI7/MM2_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI7/MM0 N_YOUT<7>_XI26/XI7/MM0_d N_Y_SEL<1>_XI26/XI7/MM0_g
+ N_VDD_XI26/XI7/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI7/MM10 N_YOUT<7>_XI26/XI7/MM10_d N_Y_SEL<0>_XI26/XI7/MM10_g
+ N_VDD_XI26/XI7/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI6/MM12 N_YOUT<6>_XI26/XI6/MM12_d N_VDD_XI26/XI6/MM12_g
+ N_VDD_XI26/XI6/MM12_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI6/MM2 N_YOUT<6>_XI26/XI6/MM2_d N_XI26/NET0116_XI26/XI6/MM2_g
+ N_VDD_XI26/XI6/MM2_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI6/MM0 N_YOUT<6>_XI26/XI6/MM0_d N_Y_SEL<1>_XI26/XI6/MM0_g
+ N_VDD_XI26/XI6/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI6/MM10 N_YOUT<6>_XI26/XI6/MM10_d N_Y_SEL<0>_XI26/XI6/MM10_g
+ N_VDD_XI26/XI6/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI5/MM12 N_YOUT<5>_XI26/XI5/MM12_d N_VDD_XI26/XI5/MM12_g
+ N_VDD_XI26/XI5/MM12_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI5/MM2 N_YOUT<5>_XI26/XI5/MM2_d N_Y_SEL<2>_XI26/XI5/MM2_g
+ N_VDD_XI26/XI5/MM2_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI5/MM0 N_YOUT<5>_XI26/XI5/MM0_d N_XI26/NET0105_XI26/XI5/MM0_g
+ N_VDD_XI26/XI5/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI5/MM10 N_YOUT<5>_XI26/XI5/MM10_d N_Y_SEL<0>_XI26/XI5/MM10_g
+ N_VDD_XI26/XI5/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI4/MM12 N_YOUT<4>_XI26/XI4/MM12_d N_VDD_XI26/XI4/MM12_g
+ N_VDD_XI26/XI4/MM12_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI4/MM2 N_YOUT<4>_XI26/XI4/MM2_d N_XI26/NET0116_XI26/XI4/MM2_g
+ N_VDD_XI26/XI4/MM2_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI4/MM0 N_YOUT<4>_XI26/XI4/MM0_d N_XI26/NET0105_XI26/XI4/MM0_g
+ N_VDD_XI26/XI4/MM0_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI4/MM10 N_YOUT<4>_XI26/XI4/MM10_d N_Y_SEL<0>_XI26/XI4/MM10_g
+ N_VDD_XI26/XI4/MM10_s N_VDD_XI26/XI7/MM12_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI26/XI10/MM10 N_XI26/NET0116_XI26/XI10/MM10_d N_Y_SEL<2>_XI26/XI10/MM10_g
+ N_VSS_XI26/XI10/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI26/XI10/MM6 N_XI26/NET0116_XI26/XI10/MM6_d N_Y_SEL<2>_XI26/XI10/MM6_g
+ N_VDD_XI26/XI10/MM6_s N_VDD_XI26/XI10/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI26/XI11/MM10 N_XI26/NET0105_XI26/XI11/MM10_d N_Y_SEL<1>_XI26/XI11/MM10_g
+ N_VSS_XI26/XI11/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI26/XI11/MM6 N_XI26/NET0105_XI26/XI11/MM6_d N_Y_SEL<1>_XI26/XI11/MM6_g
+ N_VDD_XI26/XI11/MM6_s N_VDD_XI26/XI11/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI26/XI8/MM10 N_XI26/NET0158_XI26/XI8/MM10_d N_Y_SEL<0>_XI26/XI8/MM10_g
+ N_VSS_XI26/XI8/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI26/XI8/MM6 N_XI26/NET0158_XI26/XI8/MM6_d N_Y_SEL<0>_XI26/XI8/MM6_g
+ N_VDD_XI26/XI8/MM6_s N_VDD_XI26/XI8/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13
+ AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI49/XI5/MM10 N_XI29/XI49/NET14_XI29/XI49/XI5/MM10_d
+ N_XI29/NET0150_XI29/XI49/XI5/MM10_g N_VSS_XI29/XI49/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI49/XI5/MM6 N_XI29/XI49/NET14_XI29/XI49/XI5/MM6_d
+ N_XI29/NET0150_XI29/XI49/XI5/MM6_g N_VDD_XI29/XI49/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI49/XI7/MM10 N_XI29/NET0146_XI29/XI49/XI7/MM10_d
+ N_XI29/XI49/NET14_XI29/XI49/XI7/MM10_g N_VSS_XI29/XI49/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI49/XI7/MM6 N_XI29/NET0146_XI29/XI49/XI7/MM6_d
+ N_XI29/XI49/NET14_XI29/XI49/XI7/MM6_g N_VDD_XI29/XI49/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI47/XI5/MM10 N_XI29/XI47/NET14_XI29/XI47/XI5/MM10_d
+ N_XI29/NET0130_XI29/XI47/XI5/MM10_g N_VSS_XI29/XI47/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI47/XI5/MM6 N_XI29/XI47/NET14_XI29/XI47/XI5/MM6_d
+ N_XI29/NET0130_XI29/XI47/XI5/MM6_g N_VDD_XI29/XI47/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI47/XI7/MM10 N_XI29/NET0126_XI29/XI47/XI7/MM10_d
+ N_XI29/XI47/NET14_XI29/XI47/XI7/MM10_g N_VSS_XI29/XI47/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI47/XI7/MM6 N_XI29/NET0126_XI29/XI47/XI7/MM6_d
+ N_XI29/XI47/NET14_XI29/XI47/XI7/MM6_g N_VDD_XI29/XI47/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI48/XI5/MM10 N_XI29/XI48/NET14_XI29/XI48/XI5/MM10_d
+ N_XI29/NET0126_XI29/XI48/XI5/MM10_g N_VSS_XI29/XI48/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI48/XI5/MM6 N_XI29/XI48/NET14_XI29/XI48/XI5/MM6_d
+ N_XI29/NET0126_XI29/XI48/XI5/MM6_g N_VDD_XI29/XI48/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI48/XI7/MM10 N_XI29/NET0150_XI29/XI48/XI7/MM10_d
+ N_XI29/XI48/NET14_XI29/XI48/XI7/MM10_g N_VSS_XI29/XI48/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI48/XI7/MM6 N_XI29/NET0150_XI29/XI48/XI7/MM6_d
+ N_XI29/XI48/NET14_XI29/XI48/XI7/MM6_g N_VDD_XI29/XI48/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI58/XI7/MM10 N_XI29/NET0106_XI29/XI58/XI7/MM10_d
+ N_XI29/XI58/NET14_XI29/XI58/XI7/MM10_g N_VSS_XI29/XI58/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI58/XI7/MM6 N_XI29/NET0106_XI29/XI58/XI7/MM6_d
+ N_XI29/XI58/NET14_XI29/XI58/XI7/MM6_g N_VDD_XI29/XI58/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI59/XI5/MM10 N_XI29/XI59/NET14_XI29/XI59/XI5/MM10_d
+ N_XI29/NET0106_XI29/XI59/XI5/MM10_g N_VSS_XI29/XI59/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI59/XI5/MM6 N_XI29/XI59/NET14_XI29/XI59/XI5/MM6_d
+ N_XI29/NET0106_XI29/XI59/XI5/MM6_g N_VDD_XI29/XI59/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI59/XI7/MM10 N_XI29/NET0185_XI29/XI59/XI7/MM10_d
+ N_XI29/XI59/NET14_XI29/XI59/XI7/MM10_g N_VSS_XI29/XI59/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI59/XI7/MM6 N_XI29/NET0185_XI29/XI59/XI7/MM6_d
+ N_XI29/XI59/NET14_XI29/XI59/XI7/MM6_g N_VDD_XI29/XI59/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI72/XI5/MM10 N_XI29/XI72/NET14_XI29/XI72/XI5/MM10_d
+ N_XI29/NET0185_XI29/XI72/XI5/MM10_g N_VSS_XI29/XI72/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI72/XI5/MM6 N_XI29/XI72/NET14_XI29/XI72/XI5/MM6_d
+ N_XI29/NET0185_XI29/XI72/XI5/MM6_g N_VDD_XI29/XI72/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI63/XI7/MM10 N_XI29/NET099_XI29/XI63/XI7/MM10_d
+ N_XI29/XI63/NET14_XI29/XI63/XI7/MM10_g N_VSS_XI29/XI63/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI63/XI7/MM6 N_XI29/NET099_XI29/XI63/XI7/MM6_d
+ N_XI29/XI63/NET14_XI29/XI63/XI7/MM6_g N_VDD_XI29/XI63/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI65/XI5/MM10 N_XI29/XI65/NET14_XI29/XI65/XI5/MM10_d
+ N_XI29/NET099_XI29/XI65/XI5/MM10_g N_VSS_XI29/XI65/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI65/XI5/MM6 N_XI29/XI65/NET14_XI29/XI65/XI5/MM6_d
+ N_XI29/NET099_XI29/XI65/XI5/MM6_g N_VDD_XI29/XI65/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI65/XI7/MM10 N_XI29/NET0134_XI29/XI65/XI7/MM10_d
+ N_XI29/XI65/NET14_XI29/XI65/XI7/MM10_g N_VSS_XI29/XI65/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI65/XI7/MM6 N_XI29/NET0134_XI29/XI65/XI7/MM6_d
+ N_XI29/XI65/NET14_XI29/XI65/XI7/MM6_g N_VDD_XI29/XI65/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI60/MM10 N_XI29/NET101_XI29/XI60/MM10_d N_XI29/NET0134_XI29/XI60/MM10_g
+ N_VSS_XI29/XI60/MM10_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13
+ AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI60/MM6 N_XI29/NET101_XI29/XI60/MM6_d N_XI29/NET0134_XI29/XI60/MM6_g
+ N_VDD_XI29/XI60/MM6_s N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI50/XI7/MM10 N_XI29/NET094_XI29/XI50/XI7/MM10_d
+ N_XI29/XI50/NET14_XI29/XI50/XI7/MM10_g N_VSS_XI29/XI50/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI50/XI7/MM6 N_XI29/NET094_XI29/XI50/XI7/MM6_d
+ N_XI29/XI50/NET14_XI29/XI50/XI7/MM6_g N_VDD_XI29/XI50/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI51/XI5/MM10 N_XI29/XI51/NET14_XI29/XI51/XI5/MM10_d
+ N_XI29/NET094_XI29/XI51/XI5/MM10_g N_VSS_XI29/XI51/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI51/XI5/MM6 N_XI29/XI51/NET14_XI29/XI51/XI5/MM6_d
+ N_XI29/NET094_XI29/XI51/XI5/MM6_g N_VDD_XI29/XI51/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI51/XI7/MM10 N_XI29/NET0102_XI29/XI51/XI7/MM10_d
+ N_XI29/XI51/NET14_XI29/XI51/XI7/MM10_g N_VSS_XI29/XI51/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI51/XI7/MM6 N_XI29/NET0102_XI29/XI51/XI7/MM6_d
+ N_XI29/XI51/NET14_XI29/XI51/XI7/MM6_g N_VDD_XI29/XI51/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI52/XI5/MM10 N_XI29/XI52/NET14_XI29/XI52/XI5/MM10_d
+ N_XI29/NET0102_XI29/XI52/XI5/MM10_g N_VSS_XI29/XI52/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI52/XI5/MM6 N_XI29/XI52/NET14_XI29/XI52/XI5/MM6_d
+ N_XI29/NET0102_XI29/XI52/XI5/MM6_g N_VDD_XI29/XI52/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI52/XI7/MM10 N_XI29/NET0110_XI29/XI52/XI7/MM10_d
+ N_XI29/XI52/NET14_XI29/XI52/XI7/MM10_g N_VSS_XI29/XI52/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI52/XI7/MM6 N_XI29/NET0110_XI29/XI52/XI7/MM6_d
+ N_XI29/XI52/NET14_XI29/XI52/XI7/MM6_g N_VDD_XI29/XI52/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI53/XI5/MM10 N_XI29/XI53/NET14_XI29/XI53/XI5/MM10_d
+ N_XI29/NET0110_XI29/XI53/XI5/MM10_g N_VSS_XI29/XI53/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI53/XI5/MM6 N_XI29/XI53/NET14_XI29/XI53/XI5/MM6_d
+ N_XI29/NET0110_XI29/XI53/XI5/MM6_g N_VDD_XI29/XI53/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI53/XI7/MM10 N_XI29/NET0154_XI29/XI53/XI7/MM10_d
+ N_XI29/XI53/NET14_XI29/XI53/XI7/MM10_g N_VSS_XI29/XI53/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI53/XI7/MM6 N_XI29/NET0154_XI29/XI53/XI7/MM6_d
+ N_XI29/XI53/NET14_XI29/XI53/XI7/MM6_g N_VDD_XI29/XI53/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI54/XI5/MM10 N_XI29/XI54/NET14_XI29/XI54/XI5/MM10_d
+ N_XI29/NET0154_XI29/XI54/XI5/MM10_g N_VSS_XI29/XI54/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI54/XI5/MM6 N_XI29/XI54/NET14_XI29/XI54/XI5/MM6_d
+ N_XI29/NET0154_XI29/XI54/XI5/MM6_g N_VDD_XI29/XI54/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI38/XI5/MM10 N_XI29/XI38/NET14_XI29/XI38/XI5/MM10_d
+ N_CLK_XI29/XI38/XI5/MM10_g N_VSS_XI29/XI38/XI5/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI38/XI5/MM6 N_XI29/XI38/NET14_XI29/XI38/XI5/MM6_d
+ N_CLK_XI29/XI38/XI5/MM6_g N_VDD_XI29/XI38/XI5/MM6_s N_VDD_XI29/XI50/XI5/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI38/XI7/MM10 N_XI29/NET109_XI29/XI38/XI7/MM10_d
+ N_XI29/XI38/NET14_XI29/XI38/XI7/MM10_g N_VSS_XI29/XI38/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI38/XI7/MM6 N_XI29/NET109_XI29/XI38/XI7/MM6_d
+ N_XI29/XI38/NET14_XI29/XI38/XI7/MM6_g N_VDD_XI29/XI38/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI39/XI5/MM10 N_XI29/XI39/NET14_XI29/XI39/XI5/MM10_d
+ N_XI29/NET109_XI29/XI39/XI5/MM10_g N_VSS_XI29/XI39/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI39/XI5/MM6 N_XI29/XI39/NET14_XI29/XI39/XI5/MM6_d
+ N_XI29/NET109_XI29/XI39/XI5/MM6_g N_VDD_XI29/XI39/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI39/XI7/MM10 N_XI29/NET105_XI29/XI39/XI7/MM10_d
+ N_XI29/XI39/NET14_XI29/XI39/XI7/MM10_g N_VSS_XI29/XI39/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI39/XI7/MM6 N_XI29/NET105_XI29/XI39/XI7/MM6_d
+ N_XI29/XI39/NET14_XI29/XI39/XI7/MM6_g N_VDD_XI29/XI39/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI40/XI5/MM10 N_XI29/XI40/NET14_XI29/XI40/XI5/MM10_d
+ N_XI29/NET105_XI29/XI40/XI5/MM10_g N_VSS_XI29/XI40/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI40/XI5/MM6 N_XI29/XI40/NET14_XI29/XI40/XI5/MM6_d
+ N_XI29/NET105_XI29/XI40/XI5/MM6_g N_VDD_XI29/XI40/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI40/XI7/MM10 N_XI29/NET113_XI29/XI40/XI7/MM10_d
+ N_XI29/XI40/NET14_XI29/XI40/XI7/MM10_g N_VSS_XI29/XI40/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI40/XI7/MM6 N_XI29/NET113_XI29/XI40/XI7/MM6_d
+ N_XI29/XI40/NET14_XI29/XI40/XI7/MM6_g N_VDD_XI29/XI40/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI46/XI5/MM10 N_XI29/XI46/NET14_XI29/XI46/XI5/MM10_d
+ N_XI29/NET113_XI29/XI46/XI5/MM10_g N_VSS_XI29/XI46/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI46/XI5/MM6 N_XI29/XI46/NET14_XI29/XI46/XI5/MM6_d
+ N_XI29/NET113_XI29/XI46/XI5/MM6_g N_VDD_XI29/XI46/XI5/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI46/XI7/MM10 N_XI29/NET0130_XI29/XI46/XI7/MM10_d
+ N_XI29/XI46/NET14_XI29/XI46/XI7/MM10_g N_VSS_XI29/XI46/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI46/XI7/MM6 N_XI29/NET0130_XI29/XI46/XI7/MM6_d
+ N_XI29/XI46/NET14_XI29/XI46/XI7/MM6_g N_VDD_XI29/XI46/XI7/MM6_s
+ N_VDD_XI29/XI50/XI5/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI72/XI7/MM10 N_XI29/NET0162_XI29/XI72/XI7/MM10_d
+ N_XI29/XI72/NET14_XI29/XI72/XI7/MM10_g N_VSS_XI29/XI72/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI72/XI7/MM6 N_XI29/NET0162_XI29/XI72/XI7/MM6_d
+ N_XI29/XI72/NET14_XI29/XI72/XI7/MM6_g N_VDD_XI29/XI72/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI71/XI5/MM10 N_XI29/XI71/NET14_XI29/XI71/XI5/MM10_d
+ N_XI29/NET0162_XI29/XI71/XI5/MM10_g N_VSS_XI29/XI71/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI71/XI5/MM6 N_XI29/XI71/NET14_XI29/XI71/XI5/MM6_d
+ N_XI29/NET0162_XI29/XI71/XI5/MM6_g N_VDD_XI29/XI71/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI71/XI7/MM10 N_XI29/NET0158_XI29/XI71/XI7/MM10_d
+ N_XI29/XI71/NET14_XI29/XI71/XI7/MM10_g N_VSS_XI29/XI71/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI71/XI7/MM6 N_XI29/NET0158_XI29/XI71/XI7/MM6_d
+ N_XI29/XI71/NET14_XI29/XI71/XI7/MM6_g N_VDD_XI29/XI71/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI77/XI5/MM10 N_XI29/XI77/NET14_XI29/XI77/XI5/MM10_d
+ N_XI29/NET0158_XI29/XI77/XI5/MM10_g N_VSS_XI29/XI77/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI77/XI5/MM6 N_XI29/XI77/NET14_XI29/XI77/XI5/MM6_d
+ N_XI29/NET0158_XI29/XI77/XI5/MM6_g N_VDD_XI29/XI77/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI77/XI7/MM10 N_XI29/NET0182_XI29/XI77/XI7/MM10_d
+ N_XI29/XI77/NET14_XI29/XI77/XI7/MM10_g N_VSS_XI29/XI77/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI77/XI7/MM6 N_XI29/NET0182_XI29/XI77/XI7/MM6_d
+ N_XI29/XI77/NET14_XI29/XI77/XI7/MM6_g N_VDD_XI29/XI77/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI70/XI5/MM10 N_XI29/XI70/NET14_XI29/XI70/XI5/MM10_d
+ N_XI29/NET0182_XI29/XI70/XI5/MM10_g N_VSS_XI29/XI70/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI70/XI5/MM6 N_XI29/XI70/NET14_XI29/XI70/XI5/MM6_d
+ N_XI29/NET0182_XI29/XI70/XI5/MM6_g N_VDD_XI29/XI70/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI70/XI7/MM10 N_XI29/NET097_XI29/XI70/XI7/MM10_d
+ N_XI29/XI70/NET14_XI29/XI70/XI7/MM10_g N_VSS_XI29/XI70/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI70/XI7/MM6 N_XI29/NET097_XI29/XI70/XI7/MM6_d
+ N_XI29/XI70/NET14_XI29/XI70/XI7/MM6_g N_VDD_XI29/XI70/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI69/XI5/MM10 N_XI29/XI69/NET14_XI29/XI69/XI5/MM10_d
+ N_XI29/NET097_XI29/XI69/XI5/MM10_g N_VSS_XI29/XI69/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI69/XI5/MM6 N_XI29/XI69/NET14_XI29/XI69/XI5/MM6_d
+ N_XI29/NET097_XI29/XI69/XI5/MM6_g N_VDD_XI29/XI69/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI54/XI7/MM10 N_XI29/NET0142_XI29/XI54/XI7/MM10_d
+ N_XI29/XI54/NET14_XI29/XI54/XI7/MM10_g N_VSS_XI29/XI54/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI54/XI7/MM6 N_XI29/NET0142_XI29/XI54/XI7/MM6_d
+ N_XI29/XI54/NET14_XI29/XI54/XI7/MM6_g N_VDD_XI29/XI54/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI55/XI5/MM10 N_XI29/XI55/NET14_XI29/XI55/XI5/MM10_d
+ N_XI29/NET0142_XI29/XI55/XI5/MM10_g N_VSS_XI29/XI55/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI55/XI5/MM6 N_XI29/XI55/NET14_XI29/XI55/XI5/MM6_d
+ N_XI29/NET0142_XI29/XI55/XI5/MM6_g N_VDD_XI29/XI55/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI55/XI7/MM10 N_XI29/NET098_XI29/XI55/XI7/MM10_d
+ N_XI29/XI55/NET14_XI29/XI55/XI7/MM10_g N_VSS_XI29/XI55/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI55/XI7/MM6 N_XI29/NET098_XI29/XI55/XI7/MM6_d
+ N_XI29/XI55/NET14_XI29/XI55/XI7/MM6_g N_VDD_XI29/XI55/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI56/XI5/MM10 N_XI29/XI56/NET14_XI29/XI56/XI5/MM10_d
+ N_XI29/NET098_XI29/XI56/XI5/MM10_g N_VSS_XI29/XI56/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI56/XI5/MM6 N_XI29/XI56/NET14_XI29/XI56/XI5/MM6_d
+ N_XI29/NET098_XI29/XI56/XI5/MM6_g N_VDD_XI29/XI56/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI56/XI7/MM10 N_XI29/NET0118_XI29/XI56/XI7/MM10_d
+ N_XI29/XI56/NET14_XI29/XI56/XI7/MM10_g N_VSS_XI29/XI56/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI56/XI7/MM6 N_XI29/NET0118_XI29/XI56/XI7/MM6_d
+ N_XI29/XI56/NET14_XI29/XI56/XI7/MM6_g N_VDD_XI29/XI56/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI57/XI5/MM10 N_XI29/XI57/NET14_XI29/XI57/XI5/MM10_d
+ N_XI29/NET0118_XI29/XI57/XI5/MM10_g N_VSS_XI29/XI57/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI57/XI5/MM6 N_XI29/XI57/NET14_XI29/XI57/XI5/MM6_d
+ N_XI29/NET0118_XI29/XI57/XI5/MM6_g N_VDD_XI29/XI57/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI57/XI7/MM10 N_XI29/NET0114_XI29/XI57/XI7/MM10_d
+ N_XI29/XI57/NET14_XI29/XI57/XI7/MM10_g N_VSS_XI29/XI57/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI57/XI7/MM6 N_XI29/NET0114_XI29/XI57/XI7/MM6_d
+ N_XI29/XI57/NET14_XI29/XI57/XI7/MM6_g N_VDD_XI29/XI57/XI7/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI58/XI5/MM10 N_XI29/XI58/NET14_XI29/XI58/XI5/MM10_d
+ N_XI29/NET0114_XI29/XI58/XI5/MM10_g N_VSS_XI29/XI58/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI58/XI5/MM6 N_XI29/XI58/NET14_XI29/XI58/XI5/MM6_d
+ N_XI29/NET0114_XI29/XI58/XI5/MM6_g N_VDD_XI29/XI58/XI5/MM6_s
+ N_VDD_XI29/XI58/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI69/XI7/MM10 N_XI29/NET096_XI29/XI69/XI7/MM10_d
+ N_XI29/XI69/NET14_XI29/XI69/XI7/MM10_g N_VSS_XI29/XI69/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI69/XI7/MM6 N_XI29/NET096_XI29/XI69/XI7/MM6_d
+ N_XI29/XI69/NET14_XI29/XI69/XI7/MM6_g N_VDD_XI29/XI69/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI75/XI5/MM10 N_XI29/XI75/NET14_XI29/XI75/XI5/MM10_d
+ N_XI29/NET096_XI29/XI75/XI5/MM10_g N_VSS_XI29/XI75/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI75/XI5/MM6 N_XI29/XI75/NET14_XI29/XI75/XI5/MM6_d
+ N_XI29/NET096_XI29/XI75/XI5/MM6_g N_VDD_XI29/XI75/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI75/XI7/MM10 N_XI29/NET0174_XI29/XI75/XI7/MM10_d
+ N_XI29/XI75/NET14_XI29/XI75/XI7/MM10_g N_VSS_XI29/XI75/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI75/XI7/MM6 N_XI29/NET0174_XI29/XI75/XI7/MM6_d
+ N_XI29/XI75/NET14_XI29/XI75/XI7/MM6_g N_VDD_XI29/XI75/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI74/XI5/MM10 N_XI29/XI74/NET14_XI29/XI74/XI5/MM10_d
+ N_XI29/NET0174_XI29/XI74/XI5/MM10_g N_VSS_XI29/XI74/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI74/XI5/MM6 N_XI29/XI74/NET14_XI29/XI74/XI5/MM6_d
+ N_XI29/NET0174_XI29/XI74/XI5/MM6_g N_VDD_XI29/XI74/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI74/XI7/MM10 N_XI29/NET0170_XI29/XI74/XI7/MM10_d
+ N_XI29/XI74/NET14_XI29/XI74/XI7/MM10_g N_VSS_XI29/XI74/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI74/XI7/MM6 N_XI29/NET0170_XI29/XI74/XI7/MM6_d
+ N_XI29/XI74/NET14_XI29/XI74/XI7/MM6_g N_VDD_XI29/XI74/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI61/XI5/MM10 N_XI29/XI61/NET14_XI29/XI61/XI5/MM10_d
+ N_XI29/NET0170_XI29/XI61/XI5/MM10_g N_VSS_XI29/XI61/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI61/XI5/MM6 N_XI29/XI61/NET14_XI29/XI61/XI5/MM6_d
+ N_XI29/NET0170_XI29/XI61/XI5/MM6_g N_VDD_XI29/XI61/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI61/XI7/MM10 N_XI29/NET092_XI29/XI61/XI7/MM10_d
+ N_XI29/XI61/NET14_XI29/XI61/XI7/MM10_g N_VSS_XI29/XI61/XI7/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI61/XI7/MM6 N_XI29/NET092_XI29/XI61/XI7/MM6_d
+ N_XI29/XI61/NET14_XI29/XI61/XI7/MM6_g N_VDD_XI29/XI61/XI7/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI63/XI5/MM10 N_XI29/XI63/NET14_XI29/XI63/XI5/MM10_d
+ N_XI29/NET092_XI29/XI63/XI5/MM10_g N_VSS_XI29/XI63/XI5/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI63/XI5/MM6 N_XI29/XI63/NET14_XI29/XI63/XI5/MM6_d
+ N_XI29/NET092_XI29/XI63/XI5/MM6_g N_VDD_XI29/XI63/XI5/MM6_s
+ N_VDD_XI29/XI63/XI7/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI31/MM2 N_XI29/XI31/NET18_XI29/XI31/MM2_d N_XI29/NET0145_XI29/XI31/MM2_g
+ N_XI29/XI31/NET13_XI29/XI31/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI31/XI5/MM3 N_XI29/XI31/XI5/NET5_XI29/XI31/XI5/MM3_d
+ N_CLK_XI29/XI31/XI5/MM3_g N_VSS_XI29/XI31/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI31/XI5/MM2 N_XI29/XI31/NET13_XI29/XI31/XI5/MM2_d
+ N_XI29/XI31/NET14_XI29/XI31/XI5/MM2_g N_XI29/XI31/XI5/NET5_XI29/XI31/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI31/MM4 N_XI29/XI31/NET5_XI29/XI31/MM4_d N_CLK_XI29/XI31/MM4_g
+ N_XI29/XI31/NET14_XI29/XI31/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI31/XI6/MM3 N_XI29/XI31/XI6/NET5_XI29/XI31/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI31/XI6/MM3_g N_VSS_XI29/XI31/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI31/XI6/MM2 N_XI29/XI31/NET5_XI29/XI31/XI6/MM2_d
+ N_XI29/XI31/NET1_XI29/XI31/XI6/MM2_g N_XI29/XI31/XI6/NET5_XI29/XI31/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI31/MM0 N_XI29/XI31/NET18_XI29/XI31/MM0_d N_CLK_XI29/XI31/MM0_g
+ N_XI29/XI31/NET13_XI29/XI31/MM0_s N_VDD_XI29/XI31/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI5/MM0 N_XI29/XI31/XI5/NET12_XI29/XI31/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI31/XI5/MM0_g N_VDD_XI29/XI31/XI5/MM0_s
+ N_VDD_XI29/XI31/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI5/MM1 N_XI29/XI31/NET13_XI29/XI31/XI5/MM1_d
+ N_XI29/XI31/NET14_XI29/XI31/XI5/MM1_g
+ N_XI29/XI31/XI5/NET12_XI29/XI31/XI5/MM1_s N_VDD_XI29/XI31/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI31/MM3 N_XI29/XI31/NET5_XI29/XI31/MM3_d N_XI29/NET0145_XI29/XI31/MM3_g
+ N_XI29/XI31/NET14_XI29/XI31/MM3_s N_VDD_XI29/XI31/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI6/MM0 N_XI29/XI31/XI6/NET12_XI29/XI31/XI6/MM0_d
+ N_CLK_XI29/XI31/XI6/MM0_g N_VDD_XI29/XI31/XI6/MM0_s N_VDD_XI29/XI31/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI6/MM1 N_XI29/XI31/NET5_XI29/XI31/XI6/MM1_d
+ N_XI29/XI31/NET1_XI29/XI31/XI6/MM1_g N_XI29/XI31/XI6/NET12_XI29/XI31/XI6/MM1_s
+ N_VDD_XI29/XI31/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI0/MM10 N_XI29/XI31/NET18_XI29/XI31/XI0/MM10_d
+ N_A<2>_XI29/XI31/XI0/MM10_g N_VSS_XI29/XI31/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI31/XI0/MM6 N_XI29/XI31/NET18_XI29/XI31/XI0/MM6_d
+ N_A<2>_XI29/XI31/XI0/MM6_g N_VDD_XI29/XI31/XI0/MM6_s N_VDD_XI29/XI31/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI1/MM10 N_XI29/XI31/NET14_XI29/XI31/XI1/MM10_d
+ N_XI29/XI31/NET13_XI29/XI31/XI1/MM10_g N_VSS_XI29/XI31/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI31/XI1/MM6 N_XI29/XI31/NET14_XI29/XI31/XI1/MM6_d
+ N_XI29/XI31/NET13_XI29/XI31/XI1/MM6_g N_VDD_XI29/XI31/XI1/MM6_s
+ N_VDD_XI29/XI31/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI3/MM10 N_XI29/XI31/NET1_XI29/XI31/XI3/MM10_d
+ N_XI29/XI31/NET5_XI29/XI31/XI3/MM10_g N_VSS_XI29/XI31/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI31/XI3/MM6 N_XI29/XI31/NET1_XI29/XI31/XI3/MM6_d
+ N_XI29/XI31/NET5_XI29/XI31/XI3/MM6_g N_VDD_XI29/XI31/XI3/MM6_s
+ N_VDD_XI29/XI31/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI31/XI4/MM10 N_Y_SEL<2>_XI29/XI31/XI4/MM10_d
+ N_XI29/XI31/NET1_XI29/XI31/XI4/MM10_g N_VSS_XI29/XI31/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI31/XI4/MM6 N_Y_SEL<2>_XI29/XI31/XI4/MM6_d
+ N_XI29/XI31/NET1_XI29/XI31/XI4/MM6_g N_VDD_XI29/XI31/XI4/MM6_s
+ N_VDD_XI29/XI31/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI32/MM2 N_XI29/XI32/NET18_XI29/XI32/MM2_d N_XI29/NET0145_XI29/XI32/MM2_g
+ N_XI29/XI32/NET13_XI29/XI32/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI32/XI5/MM3 N_XI29/XI32/XI5/NET5_XI29/XI32/XI5/MM3_d
+ N_CLK_XI29/XI32/XI5/MM3_g N_VSS_XI29/XI32/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI32/XI5/MM2 N_XI29/XI32/NET13_XI29/XI32/XI5/MM2_d
+ N_XI29/XI32/NET14_XI29/XI32/XI5/MM2_g N_XI29/XI32/XI5/NET5_XI29/XI32/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI32/MM4 N_XI29/XI32/NET5_XI29/XI32/MM4_d N_CLK_XI29/XI32/MM4_g
+ N_XI29/XI32/NET14_XI29/XI32/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI32/XI6/MM3 N_XI29/XI32/XI6/NET5_XI29/XI32/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI32/XI6/MM3_g N_VSS_XI29/XI32/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI32/XI6/MM2 N_XI29/XI32/NET5_XI29/XI32/XI6/MM2_d
+ N_XI29/XI32/NET1_XI29/XI32/XI6/MM2_g N_XI29/XI32/XI6/NET5_XI29/XI32/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI32/MM0 N_XI29/XI32/NET18_XI29/XI32/MM0_d N_CLK_XI29/XI32/MM0_g
+ N_XI29/XI32/NET13_XI29/XI32/MM0_s N_VDD_XI29/XI32/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI5/MM0 N_XI29/XI32/XI5/NET12_XI29/XI32/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI32/XI5/MM0_g N_VDD_XI29/XI32/XI5/MM0_s
+ N_VDD_XI29/XI32/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI5/MM1 N_XI29/XI32/NET13_XI29/XI32/XI5/MM1_d
+ N_XI29/XI32/NET14_XI29/XI32/XI5/MM1_g
+ N_XI29/XI32/XI5/NET12_XI29/XI32/XI5/MM1_s N_VDD_XI29/XI32/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI32/MM3 N_XI29/XI32/NET5_XI29/XI32/MM3_d N_XI29/NET0145_XI29/XI32/MM3_g
+ N_XI29/XI32/NET14_XI29/XI32/MM3_s N_VDD_XI29/XI32/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI6/MM0 N_XI29/XI32/XI6/NET12_XI29/XI32/XI6/MM0_d
+ N_CLK_XI29/XI32/XI6/MM0_g N_VDD_XI29/XI32/XI6/MM0_s N_VDD_XI29/XI32/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI6/MM1 N_XI29/XI32/NET5_XI29/XI32/XI6/MM1_d
+ N_XI29/XI32/NET1_XI29/XI32/XI6/MM1_g N_XI29/XI32/XI6/NET12_XI29/XI32/XI6/MM1_s
+ N_VDD_XI29/XI32/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI0/MM10 N_XI29/XI32/NET18_XI29/XI32/XI0/MM10_d
+ N_A<1>_XI29/XI32/XI0/MM10_g N_VSS_XI29/XI32/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI32/XI0/MM6 N_XI29/XI32/NET18_XI29/XI32/XI0/MM6_d
+ N_A<1>_XI29/XI32/XI0/MM6_g N_VDD_XI29/XI32/XI0/MM6_s N_VDD_XI29/XI32/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI1/MM10 N_XI29/XI32/NET14_XI29/XI32/XI1/MM10_d
+ N_XI29/XI32/NET13_XI29/XI32/XI1/MM10_g N_VSS_XI29/XI32/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI32/XI1/MM6 N_XI29/XI32/NET14_XI29/XI32/XI1/MM6_d
+ N_XI29/XI32/NET13_XI29/XI32/XI1/MM6_g N_VDD_XI29/XI32/XI1/MM6_s
+ N_VDD_XI29/XI32/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI3/MM10 N_XI29/XI32/NET1_XI29/XI32/XI3/MM10_d
+ N_XI29/XI32/NET5_XI29/XI32/XI3/MM10_g N_VSS_XI29/XI32/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI32/XI3/MM6 N_XI29/XI32/NET1_XI29/XI32/XI3/MM6_d
+ N_XI29/XI32/NET5_XI29/XI32/XI3/MM6_g N_VDD_XI29/XI32/XI3/MM6_s
+ N_VDD_XI29/XI32/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI32/XI4/MM10 N_Y_SEL<1>_XI29/XI32/XI4/MM10_d
+ N_XI29/XI32/NET1_XI29/XI32/XI4/MM10_g N_VSS_XI29/XI32/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI32/XI4/MM6 N_Y_SEL<1>_XI29/XI32/XI4/MM6_d
+ N_XI29/XI32/NET1_XI29/XI32/XI4/MM6_g N_VDD_XI29/XI32/XI4/MM6_s
+ N_VDD_XI29/XI32/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI35/MM2 N_XI29/XI35/NET18_XI29/XI35/MM2_d N_XI29/NET0145_XI29/XI35/MM2_g
+ N_XI29/XI35/NET13_XI29/XI35/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI35/XI5/MM3 N_XI29/XI35/XI5/NET5_XI29/XI35/XI5/MM3_d
+ N_CLK_XI29/XI35/XI5/MM3_g N_VSS_XI29/XI35/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI35/XI5/MM2 N_XI29/XI35/NET13_XI29/XI35/XI5/MM2_d
+ N_XI29/XI35/NET14_XI29/XI35/XI5/MM2_g N_XI29/XI35/XI5/NET5_XI29/XI35/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI35/MM4 N_XI29/XI35/NET5_XI29/XI35/MM4_d N_CLK_XI29/XI35/MM4_g
+ N_XI29/XI35/NET14_XI29/XI35/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI35/XI6/MM3 N_XI29/XI35/XI6/NET5_XI29/XI35/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI35/XI6/MM3_g N_VSS_XI29/XI35/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI35/XI6/MM2 N_XI29/XI35/NET5_XI29/XI35/XI6/MM2_d
+ N_XI29/XI35/NET1_XI29/XI35/XI6/MM2_g N_XI29/XI35/XI6/NET5_XI29/XI35/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI35/MM0 N_XI29/XI35/NET18_XI29/XI35/MM0_d N_CLK_XI29/XI35/MM0_g
+ N_XI29/XI35/NET13_XI29/XI35/MM0_s N_VDD_XI29/XI35/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI5/MM0 N_XI29/XI35/XI5/NET12_XI29/XI35/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI35/XI5/MM0_g N_VDD_XI29/XI35/XI5/MM0_s
+ N_VDD_XI29/XI35/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI5/MM1 N_XI29/XI35/NET13_XI29/XI35/XI5/MM1_d
+ N_XI29/XI35/NET14_XI29/XI35/XI5/MM1_g
+ N_XI29/XI35/XI5/NET12_XI29/XI35/XI5/MM1_s N_VDD_XI29/XI35/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI35/MM3 N_XI29/XI35/NET5_XI29/XI35/MM3_d N_XI29/NET0145_XI29/XI35/MM3_g
+ N_XI29/XI35/NET14_XI29/XI35/MM3_s N_VDD_XI29/XI35/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI6/MM0 N_XI29/XI35/XI6/NET12_XI29/XI35/XI6/MM0_d
+ N_CLK_XI29/XI35/XI6/MM0_g N_VDD_XI29/XI35/XI6/MM0_s N_VDD_XI29/XI35/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI6/MM1 N_XI29/XI35/NET5_XI29/XI35/XI6/MM1_d
+ N_XI29/XI35/NET1_XI29/XI35/XI6/MM1_g N_XI29/XI35/XI6/NET12_XI29/XI35/XI6/MM1_s
+ N_VDD_XI29/XI35/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI0/MM10 N_XI29/XI35/NET18_XI29/XI35/XI0/MM10_d
+ N_A<0>_XI29/XI35/XI0/MM10_g N_VSS_XI29/XI35/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI35/XI0/MM6 N_XI29/XI35/NET18_XI29/XI35/XI0/MM6_d
+ N_A<0>_XI29/XI35/XI0/MM6_g N_VDD_XI29/XI35/XI0/MM6_s N_VDD_XI29/XI35/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI1/MM10 N_XI29/XI35/NET14_XI29/XI35/XI1/MM10_d
+ N_XI29/XI35/NET13_XI29/XI35/XI1/MM10_g N_VSS_XI29/XI35/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI35/XI1/MM6 N_XI29/XI35/NET14_XI29/XI35/XI1/MM6_d
+ N_XI29/XI35/NET13_XI29/XI35/XI1/MM6_g N_VDD_XI29/XI35/XI1/MM6_s
+ N_VDD_XI29/XI35/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI3/MM10 N_XI29/XI35/NET1_XI29/XI35/XI3/MM10_d
+ N_XI29/XI35/NET5_XI29/XI35/XI3/MM10_g N_VSS_XI29/XI35/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI35/XI3/MM6 N_XI29/XI35/NET1_XI29/XI35/XI3/MM6_d
+ N_XI29/XI35/NET5_XI29/XI35/XI3/MM6_g N_VDD_XI29/XI35/XI3/MM6_s
+ N_VDD_XI29/XI35/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI35/XI4/MM10 N_Y_SEL<0>_XI29/XI35/XI4/MM10_d
+ N_XI29/XI35/NET1_XI29/XI35/XI4/MM10_g N_VSS_XI29/XI35/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI35/XI4/MM6 N_Y_SEL<0>_XI29/XI35/XI4/MM6_d
+ N_XI29/XI35/NET1_XI29/XI35/XI4/MM6_g N_VDD_XI29/XI35/XI4/MM6_s
+ N_VDD_XI29/XI35/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI30/MM2 N_XI29/XI30/NET18_XI29/XI30/MM2_d N_XI29/NET0145_XI29/XI30/MM2_g
+ N_XI29/XI30/NET13_XI29/XI30/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI30/XI5/MM3 N_XI29/XI30/XI5/NET5_XI29/XI30/XI5/MM3_d
+ N_CLK_XI29/XI30/XI5/MM3_g N_VSS_XI29/XI30/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI30/XI5/MM2 N_XI29/XI30/NET13_XI29/XI30/XI5/MM2_d
+ N_XI29/XI30/NET14_XI29/XI30/XI5/MM2_g N_XI29/XI30/XI5/NET5_XI29/XI30/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI30/MM4 N_XI29/XI30/NET5_XI29/XI30/MM4_d N_CLK_XI29/XI30/MM4_g
+ N_XI29/XI30/NET14_XI29/XI30/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI30/XI6/MM3 N_XI29/XI30/XI6/NET5_XI29/XI30/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI30/XI6/MM3_g N_VSS_XI29/XI30/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI30/XI6/MM2 N_XI29/XI30/NET5_XI29/XI30/XI6/MM2_d
+ N_XI29/XI30/NET1_XI29/XI30/XI6/MM2_g N_XI29/XI30/XI6/NET5_XI29/XI30/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI30/MM0 N_XI29/XI30/NET18_XI29/XI30/MM0_d N_CLK_XI29/XI30/MM0_g
+ N_XI29/XI30/NET13_XI29/XI30/MM0_s N_VDD_XI29/XI30/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI5/MM0 N_XI29/XI30/XI5/NET12_XI29/XI30/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI30/XI5/MM0_g N_VDD_XI29/XI30/XI5/MM0_s
+ N_VDD_XI29/XI30/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI5/MM1 N_XI29/XI30/NET13_XI29/XI30/XI5/MM1_d
+ N_XI29/XI30/NET14_XI29/XI30/XI5/MM1_g
+ N_XI29/XI30/XI5/NET12_XI29/XI30/XI5/MM1_s N_VDD_XI29/XI30/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI30/MM3 N_XI29/XI30/NET5_XI29/XI30/MM3_d N_XI29/NET0145_XI29/XI30/MM3_g
+ N_XI29/XI30/NET14_XI29/XI30/MM3_s N_VDD_XI29/XI30/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI6/MM0 N_XI29/XI30/XI6/NET12_XI29/XI30/XI6/MM0_d
+ N_CLK_XI29/XI30/XI6/MM0_g N_VDD_XI29/XI30/XI6/MM0_s N_VDD_XI29/XI30/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI6/MM1 N_XI29/XI30/NET5_XI29/XI30/XI6/MM1_d
+ N_XI29/XI30/NET1_XI29/XI30/XI6/MM1_g N_XI29/XI30/XI6/NET12_XI29/XI30/XI6/MM1_s
+ N_VDD_XI29/XI30/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI0/MM10 N_XI29/XI30/NET18_XI29/XI30/XI0/MM10_d
+ N_A<6>_XI29/XI30/XI0/MM10_g N_VSS_XI29/XI30/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI30/XI0/MM6 N_XI29/XI30/NET18_XI29/XI30/XI0/MM6_d
+ N_A<6>_XI29/XI30/XI0/MM6_g N_VDD_XI29/XI30/XI0/MM6_s N_VDD_XI29/XI30/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI1/MM10 N_XI29/XI30/NET14_XI29/XI30/XI1/MM10_d
+ N_XI29/XI30/NET13_XI29/XI30/XI1/MM10_g N_VSS_XI29/XI30/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI30/XI1/MM6 N_XI29/XI30/NET14_XI29/XI30/XI1/MM6_d
+ N_XI29/XI30/NET13_XI29/XI30/XI1/MM6_g N_VDD_XI29/XI30/XI1/MM6_s
+ N_VDD_XI29/XI30/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI3/MM10 N_XI29/XI30/NET1_XI29/XI30/XI3/MM10_d
+ N_XI29/XI30/NET5_XI29/XI30/XI3/MM10_g N_VSS_XI29/XI30/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI30/XI3/MM6 N_XI29/XI30/NET1_XI29/XI30/XI3/MM6_d
+ N_XI29/XI30/NET5_XI29/XI30/XI3/MM6_g N_VDD_XI29/XI30/XI3/MM6_s
+ N_VDD_XI29/XI30/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI30/XI4/MM10 N_X_SEL<3>_XI29/XI30/XI4/MM10_d
+ N_XI29/XI30/NET1_XI29/XI30/XI4/MM10_g N_VSS_XI29/XI30/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI30/XI4/MM6 N_X_SEL<3>_XI29/XI30/XI4/MM6_d
+ N_XI29/XI30/NET1_XI29/XI30/XI4/MM6_g N_VDD_XI29/XI30/XI4/MM6_s
+ N_VDD_XI29/XI30/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI28/MM2 N_XI29/XI28/NET18_XI29/XI28/MM2_d N_XI29/NET0145_XI29/XI28/MM2_g
+ N_XI29/XI28/NET13_XI29/XI28/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI28/XI5/MM3 N_XI29/XI28/XI5/NET5_XI29/XI28/XI5/MM3_d
+ N_CLK_XI29/XI28/XI5/MM3_g N_VSS_XI29/XI28/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI28/XI5/MM2 N_XI29/XI28/NET13_XI29/XI28/XI5/MM2_d
+ N_XI29/XI28/NET14_XI29/XI28/XI5/MM2_g N_XI29/XI28/XI5/NET5_XI29/XI28/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI28/MM4 N_XI29/XI28/NET5_XI29/XI28/MM4_d N_CLK_XI29/XI28/MM4_g
+ N_XI29/XI28/NET14_XI29/XI28/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI28/XI6/MM3 N_XI29/XI28/XI6/NET5_XI29/XI28/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI28/XI6/MM3_g N_VSS_XI29/XI28/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI28/XI6/MM2 N_XI29/XI28/NET5_XI29/XI28/XI6/MM2_d
+ N_XI29/XI28/NET1_XI29/XI28/XI6/MM2_g N_XI29/XI28/XI6/NET5_XI29/XI28/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI28/MM0 N_XI29/XI28/NET18_XI29/XI28/MM0_d N_CLK_XI29/XI28/MM0_g
+ N_XI29/XI28/NET13_XI29/XI28/MM0_s N_VDD_XI29/XI28/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI5/MM0 N_XI29/XI28/XI5/NET12_XI29/XI28/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI28/XI5/MM0_g N_VDD_XI29/XI28/XI5/MM0_s
+ N_VDD_XI29/XI28/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI5/MM1 N_XI29/XI28/NET13_XI29/XI28/XI5/MM1_d
+ N_XI29/XI28/NET14_XI29/XI28/XI5/MM1_g
+ N_XI29/XI28/XI5/NET12_XI29/XI28/XI5/MM1_s N_VDD_XI29/XI28/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI28/MM3 N_XI29/XI28/NET5_XI29/XI28/MM3_d N_XI29/NET0145_XI29/XI28/MM3_g
+ N_XI29/XI28/NET14_XI29/XI28/MM3_s N_VDD_XI29/XI28/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI6/MM0 N_XI29/XI28/XI6/NET12_XI29/XI28/XI6/MM0_d
+ N_CLK_XI29/XI28/XI6/MM0_g N_VDD_XI29/XI28/XI6/MM0_s N_VDD_XI29/XI28/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI6/MM1 N_XI29/XI28/NET5_XI29/XI28/XI6/MM1_d
+ N_XI29/XI28/NET1_XI29/XI28/XI6/MM1_g N_XI29/XI28/XI6/NET12_XI29/XI28/XI6/MM1_s
+ N_VDD_XI29/XI28/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI0/MM10 N_XI29/XI28/NET18_XI29/XI28/XI0/MM10_d
+ N_A<7>_XI29/XI28/XI0/MM10_g N_VSS_XI29/XI28/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI28/XI0/MM6 N_XI29/XI28/NET18_XI29/XI28/XI0/MM6_d
+ N_A<7>_XI29/XI28/XI0/MM6_g N_VDD_XI29/XI28/XI0/MM6_s N_VDD_XI29/XI28/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI1/MM10 N_XI29/XI28/NET14_XI29/XI28/XI1/MM10_d
+ N_XI29/XI28/NET13_XI29/XI28/XI1/MM10_g N_VSS_XI29/XI28/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI28/XI1/MM6 N_XI29/XI28/NET14_XI29/XI28/XI1/MM6_d
+ N_XI29/XI28/NET13_XI29/XI28/XI1/MM6_g N_VDD_XI29/XI28/XI1/MM6_s
+ N_VDD_XI29/XI28/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI3/MM10 N_XI29/XI28/NET1_XI29/XI28/XI3/MM10_d
+ N_XI29/XI28/NET5_XI29/XI28/XI3/MM10_g N_VSS_XI29/XI28/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI28/XI3/MM6 N_XI29/XI28/NET1_XI29/XI28/XI3/MM6_d
+ N_XI29/XI28/NET5_XI29/XI28/XI3/MM6_g N_VDD_XI29/XI28/XI3/MM6_s
+ N_VDD_XI29/XI28/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI28/XI4/MM10 N_X_SEL<4>_XI29/XI28/XI4/MM10_d
+ N_XI29/XI28/NET1_XI29/XI28/XI4/MM10_g N_VSS_XI29/XI28/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI28/XI4/MM6 N_X_SEL<4>_XI29/XI28/XI4/MM6_d
+ N_XI29/XI28/NET1_XI29/XI28/XI4/MM6_g N_VDD_XI29/XI28/XI4/MM6_s
+ N_VDD_XI29/XI28/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI21/MM2 N_XI29/XI21/NET18_XI29/XI21/MM2_d N_XI29/NET0145_XI29/XI21/MM2_g
+ N_XI29/XI21/NET13_XI29/XI21/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI21/XI5/MM3 N_XI29/XI21/XI5/NET5_XI29/XI21/XI5/MM3_d
+ N_CLK_XI29/XI21/XI5/MM3_g N_VSS_XI29/XI21/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI21/XI5/MM2 N_XI29/XI21/NET13_XI29/XI21/XI5/MM2_d
+ N_XI29/XI21/NET14_XI29/XI21/XI5/MM2_g N_XI29/XI21/XI5/NET5_XI29/XI21/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI21/MM4 N_XI29/XI21/NET5_XI29/XI21/MM4_d N_CLK_XI29/XI21/MM4_g
+ N_XI29/XI21/NET14_XI29/XI21/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI21/XI6/MM3 N_XI29/XI21/XI6/NET5_XI29/XI21/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI21/XI6/MM3_g N_VSS_XI29/XI21/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI21/XI6/MM2 N_XI29/XI21/NET5_XI29/XI21/XI6/MM2_d
+ N_XI29/XI21/NET1_XI29/XI21/XI6/MM2_g N_XI29/XI21/XI6/NET5_XI29/XI21/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI21/MM0 N_XI29/XI21/NET18_XI29/XI21/MM0_d N_CLK_XI29/XI21/MM0_g
+ N_XI29/XI21/NET13_XI29/XI21/MM0_s N_VDD_XI29/XI21/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI5/MM0 N_XI29/XI21/XI5/NET12_XI29/XI21/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI21/XI5/MM0_g N_VDD_XI29/XI21/XI5/MM0_s
+ N_VDD_XI29/XI21/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI5/MM1 N_XI29/XI21/NET13_XI29/XI21/XI5/MM1_d
+ N_XI29/XI21/NET14_XI29/XI21/XI5/MM1_g
+ N_XI29/XI21/XI5/NET12_XI29/XI21/XI5/MM1_s N_VDD_XI29/XI21/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI21/MM3 N_XI29/XI21/NET5_XI29/XI21/MM3_d N_XI29/NET0145_XI29/XI21/MM3_g
+ N_XI29/XI21/NET14_XI29/XI21/MM3_s N_VDD_XI29/XI21/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI6/MM0 N_XI29/XI21/XI6/NET12_XI29/XI21/XI6/MM0_d
+ N_CLK_XI29/XI21/XI6/MM0_g N_VDD_XI29/XI21/XI6/MM0_s N_VDD_XI29/XI21/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI6/MM1 N_XI29/XI21/NET5_XI29/XI21/XI6/MM1_d
+ N_XI29/XI21/NET1_XI29/XI21/XI6/MM1_g N_XI29/XI21/XI6/NET12_XI29/XI21/XI6/MM1_s
+ N_VDD_XI29/XI21/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI0/MM10 N_XI29/XI21/NET18_XI29/XI21/XI0/MM10_d
+ N_A<8>_XI29/XI21/XI0/MM10_g N_VSS_XI29/XI21/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI21/XI0/MM6 N_XI29/XI21/NET18_XI29/XI21/XI0/MM6_d
+ N_A<8>_XI29/XI21/XI0/MM6_g N_VDD_XI29/XI21/XI0/MM6_s N_VDD_XI29/XI21/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI1/MM10 N_XI29/XI21/NET14_XI29/XI21/XI1/MM10_d
+ N_XI29/XI21/NET13_XI29/XI21/XI1/MM10_g N_VSS_XI29/XI21/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI21/XI1/MM6 N_XI29/XI21/NET14_XI29/XI21/XI1/MM6_d
+ N_XI29/XI21/NET13_XI29/XI21/XI1/MM6_g N_VDD_XI29/XI21/XI1/MM6_s
+ N_VDD_XI29/XI21/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI3/MM10 N_XI29/XI21/NET1_XI29/XI21/XI3/MM10_d
+ N_XI29/XI21/NET5_XI29/XI21/XI3/MM10_g N_VSS_XI29/XI21/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI21/XI3/MM6 N_XI29/XI21/NET1_XI29/XI21/XI3/MM6_d
+ N_XI29/XI21/NET5_XI29/XI21/XI3/MM6_g N_VDD_XI29/XI21/XI3/MM6_s
+ N_VDD_XI29/XI21/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI21/XI4/MM10 N_X_SEL<5>_XI29/XI21/XI4/MM10_d
+ N_XI29/XI21/NET1_XI29/XI21/XI4/MM10_g N_VSS_XI29/XI21/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI21/XI4/MM6 N_X_SEL<5>_XI29/XI21/XI4/MM6_d
+ N_XI29/XI21/NET1_XI29/XI21/XI4/MM6_g N_VDD_XI29/XI21/XI4/MM6_s
+ N_VDD_XI29/XI21/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI33/MM2 N_XI29/XI33/NET18_XI29/XI33/MM2_d N_XI29/NET0145_XI29/XI33/MM2_g
+ N_XI29/XI33/NET13_XI29/XI33/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI33/XI5/MM3 N_XI29/XI33/XI5/NET5_XI29/XI33/XI5/MM3_d
+ N_CLK_XI29/XI33/XI5/MM3_g N_VSS_XI29/XI33/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI33/XI5/MM2 N_XI29/XI33/NET13_XI29/XI33/XI5/MM2_d
+ N_XI29/XI33/NET14_XI29/XI33/XI5/MM2_g N_XI29/XI33/XI5/NET5_XI29/XI33/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI33/MM4 N_XI29/XI33/NET5_XI29/XI33/MM4_d N_CLK_XI29/XI33/MM4_g
+ N_XI29/XI33/NET14_XI29/XI33/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI33/XI6/MM3 N_XI29/XI33/XI6/NET5_XI29/XI33/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI33/XI6/MM3_g N_VSS_XI29/XI33/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI33/XI6/MM2 N_XI29/XI33/NET5_XI29/XI33/XI6/MM2_d
+ N_XI29/XI33/NET1_XI29/XI33/XI6/MM2_g N_XI29/XI33/XI6/NET5_XI29/XI33/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI33/MM0 N_XI29/XI33/NET18_XI29/XI33/MM0_d N_CLK_XI29/XI33/MM0_g
+ N_XI29/XI33/NET13_XI29/XI33/MM0_s N_VDD_XI29/XI33/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI5/MM0 N_XI29/XI33/XI5/NET12_XI29/XI33/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI33/XI5/MM0_g N_VDD_XI29/XI33/XI5/MM0_s
+ N_VDD_XI29/XI33/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI5/MM1 N_XI29/XI33/NET13_XI29/XI33/XI5/MM1_d
+ N_XI29/XI33/NET14_XI29/XI33/XI5/MM1_g
+ N_XI29/XI33/XI5/NET12_XI29/XI33/XI5/MM1_s N_VDD_XI29/XI33/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI33/MM3 N_XI29/XI33/NET5_XI29/XI33/MM3_d N_XI29/NET0145_XI29/XI33/MM3_g
+ N_XI29/XI33/NET14_XI29/XI33/MM3_s N_VDD_XI29/XI33/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI6/MM0 N_XI29/XI33/XI6/NET12_XI29/XI33/XI6/MM0_d
+ N_CLK_XI29/XI33/XI6/MM0_g N_VDD_XI29/XI33/XI6/MM0_s N_VDD_XI29/XI33/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI6/MM1 N_XI29/XI33/NET5_XI29/XI33/XI6/MM1_d
+ N_XI29/XI33/NET1_XI29/XI33/XI6/MM1_g N_XI29/XI33/XI6/NET12_XI29/XI33/XI6/MM1_s
+ N_VDD_XI29/XI33/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI0/MM10 N_XI29/XI33/NET18_XI29/XI33/XI0/MM10_d
+ N_A<3>_XI29/XI33/XI0/MM10_g N_VSS_XI29/XI33/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI33/XI0/MM6 N_XI29/XI33/NET18_XI29/XI33/XI0/MM6_d
+ N_A<3>_XI29/XI33/XI0/MM6_g N_VDD_XI29/XI33/XI0/MM6_s N_VDD_XI29/XI33/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI1/MM10 N_XI29/XI33/NET14_XI29/XI33/XI1/MM10_d
+ N_XI29/XI33/NET13_XI29/XI33/XI1/MM10_g N_VSS_XI29/XI33/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI33/XI1/MM6 N_XI29/XI33/NET14_XI29/XI33/XI1/MM6_d
+ N_XI29/XI33/NET13_XI29/XI33/XI1/MM6_g N_VDD_XI29/XI33/XI1/MM6_s
+ N_VDD_XI29/XI33/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI3/MM10 N_XI29/XI33/NET1_XI29/XI33/XI3/MM10_d
+ N_XI29/XI33/NET5_XI29/XI33/XI3/MM10_g N_VSS_XI29/XI33/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI33/XI3/MM6 N_XI29/XI33/NET1_XI29/XI33/XI3/MM6_d
+ N_XI29/XI33/NET5_XI29/XI33/XI3/MM6_g N_VDD_XI29/XI33/XI3/MM6_s
+ N_VDD_XI29/XI33/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI33/XI4/MM10 N_X_SEL<0>_XI29/XI33/XI4/MM10_d
+ N_XI29/XI33/NET1_XI29/XI33/XI4/MM10_g N_VSS_XI29/XI33/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI33/XI4/MM6 N_X_SEL<0>_XI29/XI33/XI4/MM6_d
+ N_XI29/XI33/NET1_XI29/XI33/XI4/MM6_g N_VDD_XI29/XI33/XI4/MM6_s
+ N_VDD_XI29/XI33/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI34/MM2 N_XI29/XI34/NET18_XI29/XI34/MM2_d N_XI29/NET0145_XI29/XI34/MM2_g
+ N_XI29/XI34/NET13_XI29/XI34/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI34/XI5/MM3 N_XI29/XI34/XI5/NET5_XI29/XI34/XI5/MM3_d
+ N_CLK_XI29/XI34/XI5/MM3_g N_VSS_XI29/XI34/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI34/XI5/MM2 N_XI29/XI34/NET13_XI29/XI34/XI5/MM2_d
+ N_XI29/XI34/NET14_XI29/XI34/XI5/MM2_g N_XI29/XI34/XI5/NET5_XI29/XI34/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI34/MM4 N_XI29/XI34/NET5_XI29/XI34/MM4_d N_CLK_XI29/XI34/MM4_g
+ N_XI29/XI34/NET14_XI29/XI34/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI34/XI6/MM3 N_XI29/XI34/XI6/NET5_XI29/XI34/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI34/XI6/MM3_g N_VSS_XI29/XI34/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI34/XI6/MM2 N_XI29/XI34/NET5_XI29/XI34/XI6/MM2_d
+ N_XI29/XI34/NET1_XI29/XI34/XI6/MM2_g N_XI29/XI34/XI6/NET5_XI29/XI34/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI34/MM0 N_XI29/XI34/NET18_XI29/XI34/MM0_d N_CLK_XI29/XI34/MM0_g
+ N_XI29/XI34/NET13_XI29/XI34/MM0_s N_VDD_XI29/XI34/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI5/MM0 N_XI29/XI34/XI5/NET12_XI29/XI34/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI34/XI5/MM0_g N_VDD_XI29/XI34/XI5/MM0_s
+ N_VDD_XI29/XI34/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI5/MM1 N_XI29/XI34/NET13_XI29/XI34/XI5/MM1_d
+ N_XI29/XI34/NET14_XI29/XI34/XI5/MM1_g
+ N_XI29/XI34/XI5/NET12_XI29/XI34/XI5/MM1_s N_VDD_XI29/XI34/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI34/MM3 N_XI29/XI34/NET5_XI29/XI34/MM3_d N_XI29/NET0145_XI29/XI34/MM3_g
+ N_XI29/XI34/NET14_XI29/XI34/MM3_s N_VDD_XI29/XI34/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI6/MM0 N_XI29/XI34/XI6/NET12_XI29/XI34/XI6/MM0_d
+ N_CLK_XI29/XI34/XI6/MM0_g N_VDD_XI29/XI34/XI6/MM0_s N_VDD_XI29/XI34/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI6/MM1 N_XI29/XI34/NET5_XI29/XI34/XI6/MM1_d
+ N_XI29/XI34/NET1_XI29/XI34/XI6/MM1_g N_XI29/XI34/XI6/NET12_XI29/XI34/XI6/MM1_s
+ N_VDD_XI29/XI34/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI0/MM10 N_XI29/XI34/NET18_XI29/XI34/XI0/MM10_d
+ N_A<4>_XI29/XI34/XI0/MM10_g N_VSS_XI29/XI34/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI34/XI0/MM6 N_XI29/XI34/NET18_XI29/XI34/XI0/MM6_d
+ N_A<4>_XI29/XI34/XI0/MM6_g N_VDD_XI29/XI34/XI0/MM6_s N_VDD_XI29/XI34/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI1/MM10 N_XI29/XI34/NET14_XI29/XI34/XI1/MM10_d
+ N_XI29/XI34/NET13_XI29/XI34/XI1/MM10_g N_VSS_XI29/XI34/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI34/XI1/MM6 N_XI29/XI34/NET14_XI29/XI34/XI1/MM6_d
+ N_XI29/XI34/NET13_XI29/XI34/XI1/MM6_g N_VDD_XI29/XI34/XI1/MM6_s
+ N_VDD_XI29/XI34/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI3/MM10 N_XI29/XI34/NET1_XI29/XI34/XI3/MM10_d
+ N_XI29/XI34/NET5_XI29/XI34/XI3/MM10_g N_VSS_XI29/XI34/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI34/XI3/MM6 N_XI29/XI34/NET1_XI29/XI34/XI3/MM6_d
+ N_XI29/XI34/NET5_XI29/XI34/XI3/MM6_g N_VDD_XI29/XI34/XI3/MM6_s
+ N_VDD_XI29/XI34/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI34/XI4/MM10 N_X_SEL<1>_XI29/XI34/XI4/MM10_d
+ N_XI29/XI34/NET1_XI29/XI34/XI4/MM10_g N_VSS_XI29/XI34/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI34/XI4/MM6 N_X_SEL<1>_XI29/XI34/XI4/MM6_d
+ N_XI29/XI34/NET1_XI29/XI34/XI4/MM6_g N_VDD_XI29/XI34/XI4/MM6_s
+ N_VDD_XI29/XI34/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI29/MM2 N_XI29/XI29/NET18_XI29/XI29/MM2_d N_XI29/NET0145_XI29/XI29/MM2_g
+ N_XI29/XI29/NET13_XI29/XI29/MM2_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI29/XI5/MM3 N_XI29/XI29/XI5/NET5_XI29/XI29/XI5/MM3_d
+ N_CLK_XI29/XI29/XI5/MM3_g N_VSS_XI29/XI29/XI5/MM3_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI29/XI5/MM2 N_XI29/XI29/NET13_XI29/XI29/XI5/MM2_d
+ N_XI29/XI29/NET14_XI29/XI29/XI5/MM2_g N_XI29/XI29/XI5/NET5_XI29/XI29/XI5/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI29/MM4 N_XI29/XI29/NET5_XI29/XI29/MM4_d N_CLK_XI29/XI29/MM4_g
+ N_XI29/XI29/NET14_XI29/XI29/MM4_s N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI29/XI6/MM3 N_XI29/XI29/XI6/NET5_XI29/XI29/XI6/MM3_d
+ N_XI29/NET0145_XI29/XI29/XI6/MM3_g N_VSS_XI29/XI29/XI6/MM3_s N_VSS_XI27/MM16_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI29/XI6/MM2 N_XI29/XI29/NET5_XI29/XI29/XI6/MM2_d
+ N_XI29/XI29/NET1_XI29/XI29/XI6/MM2_g N_XI29/XI29/XI6/NET5_XI29/XI29/XI6/MM2_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI29/MM0 N_XI29/XI29/NET18_XI29/XI29/MM0_d N_CLK_XI29/XI29/MM0_g
+ N_XI29/XI29/NET13_XI29/XI29/MM0_s N_VDD_XI29/XI29/MM0_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI5/MM0 N_XI29/XI29/XI5/NET12_XI29/XI29/XI5/MM0_d
+ N_XI29/NET0145_XI29/XI29/XI5/MM0_g N_VDD_XI29/XI29/XI5/MM0_s
+ N_VDD_XI29/XI29/XI5/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI5/MM1 N_XI29/XI29/NET13_XI29/XI29/XI5/MM1_d
+ N_XI29/XI29/NET14_XI29/XI29/XI5/MM1_g
+ N_XI29/XI29/XI5/NET12_XI29/XI29/XI5/MM1_s N_VDD_XI29/XI29/XI5/MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI29/MM3 N_XI29/XI29/NET5_XI29/XI29/MM3_d N_XI29/NET0145_XI29/XI29/MM3_g
+ N_XI29/XI29/NET14_XI29/XI29/MM3_s N_VDD_XI29/XI29/MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI6/MM0 N_XI29/XI29/XI6/NET12_XI29/XI29/XI6/MM0_d
+ N_CLK_XI29/XI29/XI6/MM0_g N_VDD_XI29/XI29/XI6/MM0_s N_VDD_XI29/XI29/XI6/MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI6/MM1 N_XI29/XI29/NET5_XI29/XI29/XI6/MM1_d
+ N_XI29/XI29/NET1_XI29/XI29/XI6/MM1_g N_XI29/XI29/XI6/NET12_XI29/XI29/XI6/MM1_s
+ N_VDD_XI29/XI29/XI6/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI0/MM10 N_XI29/XI29/NET18_XI29/XI29/XI0/MM10_d
+ N_A<5>_XI29/XI29/XI0/MM10_g N_VSS_XI29/XI29/XI0/MM10_s N_VSS_XI27/MM16_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06
mXI29/XI29/XI0/MM6 N_XI29/XI29/NET18_XI29/XI29/XI0/MM6_d
+ N_A<5>_XI29/XI29/XI0/MM6_g N_VDD_XI29/XI29/XI0/MM6_s N_VDD_XI29/XI29/XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI1/MM10 N_XI29/XI29/NET14_XI29/XI29/XI1/MM10_d
+ N_XI29/XI29/NET13_XI29/XI29/XI1/MM10_g N_VSS_XI29/XI29/XI1/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI29/XI1/MM6 N_XI29/XI29/NET14_XI29/XI29/XI1/MM6_d
+ N_XI29/XI29/NET13_XI29/XI29/XI1/MM6_g N_VDD_XI29/XI29/XI1/MM6_s
+ N_VDD_XI29/XI29/XI1/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI3/MM10 N_XI29/XI29/NET1_XI29/XI29/XI3/MM10_d
+ N_XI29/XI29/NET5_XI29/XI29/XI3/MM10_g N_VSS_XI29/XI29/XI3/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI29/XI3/MM6 N_XI29/XI29/NET1_XI29/XI29/XI3/MM6_d
+ N_XI29/XI29/NET5_XI29/XI29/XI3/MM6_g N_VDD_XI29/XI29/XI3/MM6_s
+ N_VDD_XI29/XI29/XI3/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
mXI29/XI29/XI4/MM10 N_X_SEL<2>_XI29/XI29/XI4/MM10_d
+ N_XI29/XI29/NET1_XI29/XI29/XI4/MM10_g N_VSS_XI29/XI29/XI4/MM10_s
+ N_VSS_XI27/MM16_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06
+ PS=1.52e-06
mXI29/XI29/XI4/MM6 N_X_SEL<2>_XI29/XI29/XI4/MM6_d
+ N_XI29/XI29/NET1_XI29/XI29/XI4/MM6_g N_VDD_XI29/XI29/XI4/MM6_s
+ N_VDD_XI29/XI29/XI4/MM6_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13
+ PD=2.52e-06 PS=2.52e-06
c_1 XI10/NET3768 0 0.136315f
c_2 XI10/NET5060 0 0.136314f
c_3 XI10/NET3860 0 0.136314f
c_4 XI10/NET5096 0 0.136314f
c_5 XI10/NET4104 0 0.136314f
c_6 XI10/NET3500 0 0.136314f
c_7 XI10/NET4032 0 0.136314f
c_8 XI10/NET4232 0 0.136314f
c_9 XI10/NET4572 0 0.136314f
c_10 XI10/NET4792 0 0.136314f
c_11 XI10/NET4500 0 0.136314f
c_12 XI10/NET4896 0 0.136314f
c_13 XI10/NET5456 0 0.136314f
c_14 XI10/NET5236 0 0.136314f
c_15 XI10/NET4328 0 0.136314f
c_16 XI10/NET5484 0 0.136314f
c_17 XI10/NET2136 0 0.136314f
c_18 XI10/NET2356 0 0.136314f
c_19 XI10/NET2064 0 0.136314f
c_20 XI10/NET2460 0 0.136314f
c_21 XI10/NET2844 0 0.136314f
c_22 XI10/NET02641 0 0.136314f
c_23 XI10/NET2916 0 0.136314f
c_24 XI10/NET2848 0 0.136314f
c_25 XI10/NET5632 0 0.136314f
c_26 XI10/NET1872 0 0.136314f
c_27 XI10/NET5560 0 0.136314f
c_28 XI10/NET5764 0 0.136314f
c_29 XI10/NET3088 0 0.136314f
c_30 XI10/NET3308 0 0.136314f
c_31 XI10/NET1992 0 0.136314f
c_32 XI10/NET5804 0 0.136314f
c_33 XI10/NET3720 0 0.18051f
c_34 XI10/NET5092 0 0.176433f
c_35 XI10/NET4936 0 0.176433f
c_36 XI10/NET4968 0 0.176433f
c_37 XI10/NET4172 0 0.176433f
c_38 XI10/NET4260 0 0.176433f
c_39 XI10/NET3968 0 0.176433f
c_40 XI10/NET4112 0 0.176433f
c_41 XI10/NET4640 0 0.18066f
c_42 XI10/NET4728 0 0.176433f
c_43 XI10/NET4876 0 0.176433f
c_44 XI10/NET4888 0 0.176433f
c_45 XI10/NET5388 0 0.176433f
c_46 XI10/NET5320 0 0.176433f
c_47 XI10/NET5488 0 0.176433f
c_48 XI10/NET5476 0 0.176433f
c_49 XI10/NET2204 0 0.18066f
c_50 XI10/NET2292 0 0.176433f
c_51 XI10/NET3016 0 0.176433f
c_52 XI10/NET2452 0 0.176433f
c_53 XI10/NET2776 0 0.176433f
c_54 XI10/NET2708 0 0.176433f
c_55 XI10/NET2964 0 0.176433f
c_56 XI10/NET2856 0 0.176433f
c_57 XI10/NET5700 0 0.18066f
c_58 XI10/NET5792 0 0.176433f
c_59 XI10/NET5496 0 0.176433f
c_60 XI10/NET5640 0 0.176433f
c_61 XI10/NET3156 0 0.176433f
c_62 XI10/NET3244 0 0.176433f
c_63 XI10/NET3436 0 0.176433f
c_64 XI10/NET5796 0 0.176433f
c_65 XI10/NET3732 0 0.176433f
c_66 XI10/NET5056 0 0.176433f
c_67 XI10/NET3856 0 0.176433f
c_68 XI10/NET5000 0 0.176433f
c_69 XI10/NET4100 0 0.176433f
c_70 XI10/NET3492 0 0.176433f
c_71 XI10/NET4024 0 0.176433f
c_72 XI10/NET4192 0 0.176433f
c_73 XI10/NET4568 0 0.176433f
c_74 XI10/NET4784 0 0.176433f
c_75 XI10/NET4492 0 0.176433f
c_76 XI10/NET4880 0 0.176433f
c_77 XI10/NET5448 0 0.176433f
c_78 XI10/NET5232 0 0.176433f
c_79 XI10/NET4324 0 0.176433f
c_80 XI10/NET5468 0 0.176433f
c_81 XI10/NET2132 0 0.176433f
c_82 XI10/NET2348 0 0.176433f
c_83 XI10/NET2056 0 0.176433f
c_84 XI10/NET2444 0 0.176433f
c_85 XI10/NET2836 0 0.176433f
c_86 XI10/NET02644 0 0.176433f
c_87 XI10/NET2912 0 0.176433f
c_88 XI10/NET2700 0 0.176433f
c_89 XI10/NET5628 0 0.176433f
c_90 XI10/NET1868 0 0.176433f
c_91 XI10/NET5552 0 0.176433f
c_92 XI10/NET5724 0 0.176433f
c_93 XI10/NET3084 0 0.176433f
c_94 XI10/NET3300 0 0.176433f
c_95 XI10/NET1984 0 0.176433f
c_96 XI10/NET4264 0 0.176433f
c_97 XI10/NET3712 0 0.18051f
c_98 XI10/NET5080 0 0.176433f
c_99 XI10/NET4920 0 0.176433f
c_100 XI10/NET4964 0 0.176433f
c_101 XI10/NET4168 0 0.176433f
c_102 XI10/NET4248 0 0.176433f
c_103 XI10/NET3960 0 0.176433f
c_104 XI10/NET4036 0 0.176433f
c_105 XI10/NET4636 0 0.18066f
c_106 XI10/NET4716 0 0.176433f
c_107 XI10/NET4860 0 0.176433f
c_108 XI10/NET4864 0 0.176433f
c_109 XI10/NET5380 0 0.176433f
c_110 XI10/NET5316 0 0.176433f
c_111 XI10/NET5112 0 0.176433f
c_112 XI10/NET5392 0 0.176433f
c_113 XI10/NET2200 0 0.18066f
c_114 XI10/NET2280 0 0.176433f
c_115 XI10/NET3004 0 0.176433f
c_116 XI10/NET2428 0 0.176433f
c_117 XI10/NET2768 0 0.176433f
c_118 XI10/NET2704 0 0.176433f
c_119 XI10/NET2960 0 0.176433f
c_120 XI10/NET2780 0 0.176433f
c_121 XI10/NET5696 0 0.18066f
c_122 XI10/NET5780 0 0.176433f
c_123 XI10/NET3432 0 0.176433f
c_124 XI10/NET5564 0 0.176433f
c_125 XI10/NET3152 0 0.176433f
c_126 XI10/NET3232 0 0.176433f
c_127 XI10/NET3416 0 0.176433f
c_128 XI10/NET3420 0 0.176433f
c_129 XI10/NET3752 0 0.176433f
c_130 XI10/NET5044 0 0.176433f
c_131 XI10/NET3844 0 0.176433f
c_132 XI10/NET4988 0 0.176433f
c_133 XI10/NET4088 0 0.176433f
c_134 XI10/NET3480 0 0.176433f
c_135 XI10/NET4012 0 0.176433f
c_136 XI10/NET4044 0 0.176433f
c_137 XI10/NET4556 0 0.176433f
c_138 XI10/NET4772 0 0.176433f
c_139 XI10/NET4480 0 0.176433f
c_140 XI10/NET4812 0 0.176433f
c_141 XI10/NET5436 0 0.176433f
c_142 XI10/NET5220 0 0.176433f
c_143 XI10/NET4312 0 0.176433f
c_144 XI10/NET5460 0 0.176433f
c_145 XI10/NET2120 0 0.176433f
c_146 XI10/NET2336 0 0.176433f
c_147 XI10/NET2044 0 0.176433f
c_148 XI10/NET2376 0 0.176433f
c_149 XI10/NET2824 0 0.176433f
c_150 XI10/NET02632 0 0.176433f
c_151 XI10/NET2900 0 0.176433f
c_152 XI10/NET2660 0 0.176433f
c_153 XI10/NET5616 0 0.176433f
c_154 XI10/NET1856 0 0.176433f
c_155 XI10/NET5540 0 0.176433f
c_156 XI10/NET5572 0 0.176433f
c_157 XI10/NET3072 0 0.176433f
c_158 XI10/NET3288 0 0.176433f
c_159 XI10/NET1972 0 0.176433f
c_160 XI10/NET3360 0 0.176433f
c_161 XI10/NET3700 0 0.18051f
c_162 XI10/NET5068 0 0.176433f
c_163 XI10/NET3908 0 0.176433f
c_164 XI10/NET4952 0 0.176433f
c_165 XI10/NET4156 0 0.176433f
c_166 XI10/NET4236 0 0.176433f
c_167 XI10/NET3948 0 0.176433f
c_168 XI10/NET3596 0 0.176433f
c_169 XI10/NET4624 0 0.18066f
c_170 XI10/NET4704 0 0.176433f
c_171 XI10/NET4436 0 0.176433f
c_172 XI10/NET4848 0 0.176433f
c_173 XI10/NET5368 0 0.176433f
c_174 XI10/NET5300 0 0.176433f
c_175 XI10/NET4376 0 0.176433f
c_176 XI10/NET5144 0 0.176433f
c_177 XI10/NET2188 0 0.18066f
c_178 XI10/NET2268 0 0.176433f
c_179 XI10/NET3000 0 0.176433f
c_180 XI10/NET2412 0 0.176433f
c_181 XI10/NET2756 0 0.176433f
c_182 XI10/NET2688 0 0.176433f
c_183 XI10/NET2948 0 0.176433f
c_184 XI10/NET2532 0 0.176433f
c_185 XI10/NET5684 0 0.18066f
c_186 XI10/NET5768 0 0.176433f
c_187 XI10/NET3356 0 0.176433f
c_188 XI10/NET1780 0 0.176433f
c_189 XI10/NET3140 0 0.176433f
c_190 XI10/NET3220 0 0.176433f
c_191 XI10/NET1928 0 0.176433f
c_192 XI10/NET3404 0 0.176433f
c_193 XI10/NET3780 0 0.176433f
c_194 XI10/NET5040 0 0.176433f
c_195 XI10/NET3840 0 0.176433f
c_196 XI10/NET4984 0 0.176433f
c_197 XI10/NET4084 0 0.176433f
c_198 XI10/NET3476 0 0.176433f
c_199 XI10/NET4008 0 0.176433f
c_200 XI10/NET3604 0 0.176433f
c_201 XI10/NET4552 0 0.176433f
c_202 XI10/NET4768 0 0.176433f
c_203 XI10/NET4476 0 0.176433f
c_204 XI10/NET4808 0 0.176433f
c_205 XI10/NET5432 0 0.176433f
c_206 XI10/NET5216 0 0.176433f
c_207 XI10/NET4308 0 0.176433f
c_208 XI10/NET5312 0 0.176433f
c_209 XI10/NET2116 0 0.176433f
c_210 XI10/NET2332 0 0.176433f
c_211 XI10/NET2040 0 0.176433f
c_212 XI10/NET2372 0 0.176433f
c_213 XI10/NET2820 0 0.176433f
c_214 XI10/NET02628 0 0.176433f
c_215 XI10/NET2896 0 0.176433f
c_216 XI10/NET2564 0 0.176433f
c_217 XI10/NET5612 0 0.176433f
c_218 XI10/NET1852 0 0.176433f
c_219 XI10/NET5536 0 0.176433f
c_220 XI10/NET1812 0 0.176433f
c_221 XI10/NET3068 0 0.176433f
c_222 XI10/NET3284 0 0.176433f
c_223 XI10/NET1968 0 0.176433f
c_224 XI10/NET3348 0 0.176433f
c_225 XI10/NET3696 0 0.18051f
c_226 XI10/NET3652 0 0.176433f
c_227 XI10/NET3904 0 0.176433f
c_228 XI10/NET4948 0 0.176433f
c_229 XI10/NET4152 0 0.176433f
c_230 XI10/NET4228 0 0.176433f
c_231 XI10/NET3944 0 0.176433f
c_232 XI10/NET3572 0 0.176433f
c_233 XI10/NET4620 0 0.18066f
c_234 XI10/NET4696 0 0.176433f
c_235 XI10/NET4428 0 0.176433f
c_236 XI10/NET4844 0 0.176433f
c_237 XI10/NET5364 0 0.176433f
c_238 XI10/NET5292 0 0.176433f
c_239 XI10/NET4372 0 0.176433f
c_240 XI10/NET5140 0 0.176433f
c_241 XI10/NET2184 0 0.18066f
c_242 XI10/NET2260 0 0.176433f
c_243 XI10/NET2988 0 0.176433f
c_244 XI10/NET2408 0 0.176433f
c_245 XI10/NET2752 0 0.176433f
c_246 XI10/NET2680 0 0.176433f
c_247 XI10/NET2944 0 0.176433f
c_248 XI10/NET2528 0 0.176433f
c_249 XI10/NET5680 0 0.18066f
c_250 XI10/NET5760 0 0.176433f
c_251 XI10/NET3352 0 0.176433f
c_252 XI10/NET1776 0 0.176433f
c_253 XI10/NET3136 0 0.176433f
c_254 XI10/NET3212 0 0.176433f
c_255 XI10/NET1920 0 0.176433f
c_256 XI10/NET3400 0 0.176433f
c_257 XI10/NET3748 0 0.176433f
c_258 XI10/NET5028 0 0.176433f
c_259 XI10/NET3828 0 0.176433f
c_260 XI10/NET4916 0 0.176433f
c_261 XI10/NET4072 0 0.176433f
c_262 XI10/NET3464 0 0.176433f
c_263 XI10/NET3996 0 0.176433f
c_264 XI10/NET3588 0 0.176433f
c_265 XI10/NET4540 0 0.176433f
c_266 XI10/NET4756 0 0.176433f
c_267 XI10/NET4464 0 0.176433f
c_268 XI10/NET4796 0 0.176433f
c_269 XI10/NET5420 0 0.176433f
c_270 XI10/NET5204 0 0.176433f
c_271 XI10/NET4296 0 0.176433f
c_272 XI10/NET5272 0 0.176433f
c_273 XI10/NET2104 0 0.176433f
c_274 XI10/NET2320 0 0.176433f
c_275 XI10/NET2028 0 0.176433f
c_276 XI10/NET2360 0 0.176433f
c_277 XI10/NET2808 0 0.176433f
c_278 XI10/NET02616 0 0.176433f
c_279 XI10/NET2884 0 0.176433f
c_280 XI10/NET2552 0 0.176433f
c_281 XI10/NET5600 0 0.176433f
c_282 XI10/NET1840 0 0.176433f
c_283 XI10/NET5524 0 0.176433f
c_284 XI10/NET1800 0 0.176433f
c_285 XI10/NET3056 0 0.176433f
c_286 XI10/NET3272 0 0.176433f
c_287 XI10/NET1956 0 0.176433f
c_288 XI10/NET3336 0 0.176433f
c_289 XI10/NET3684 0 0.18051f
c_290 XI10/NET3648 0 0.176433f
c_291 XI10/NET3892 0 0.176433f
c_292 XI10/NET4932 0 0.176433f
c_293 XI10/NET4140 0 0.176433f
c_294 XI10/NET4212 0 0.176433f
c_295 XI10/NET3932 0 0.176433f
c_296 XI10/NET3556 0 0.176433f
c_297 XI10/NET4608 0 0.18066f
c_298 XI10/NET4680 0 0.176433f
c_299 XI10/NET4416 0 0.176433f
c_300 XI10/NET4832 0 0.176433f
c_301 XI10/NET5352 0 0.176433f
c_302 XI10/NET5276 0 0.176433f
c_303 XI10/NET4360 0 0.176433f
c_304 XI10/NET5128 0 0.176433f
c_305 XI10/NET2172 0 0.18066f
c_306 XI10/NET2244 0 0.176433f
c_307 XI10/NET2984 0 0.176433f
c_308 XI10/NET2396 0 0.176433f
c_309 XI10/NET2740 0 0.176433f
c_310 XI10/NET2664 0 0.176433f
c_311 XI10/NET2932 0 0.176433f
c_312 XI10/NET2516 0 0.176433f
c_313 XI10/NET5668 0 0.18066f
c_314 XI10/NET5744 0 0.176433f
c_315 XI10/NET3324 0 0.176433f
c_316 XI10/NET1764 0 0.176433f
c_317 XI10/NET3124 0 0.176433f
c_318 XI10/NET3196 0 0.176433f
c_319 XI10/NET1908 0 0.176433f
c_320 XI10/NET3388 0 0.176433f
c_321 XI10/NET3764 0 0.176433f
c_322 XI10/NET5024 0 0.176433f
c_323 XI10/NET3824 0 0.176433f
c_324 XI10/NET4900 0 0.176433f
c_325 XI10/NET4068 0 0.176433f
c_326 XI10/NET3460 0 0.176433f
c_327 XI10/NET3992 0 0.176433f
c_328 XI10/NET3520 0 0.176433f
c_329 XI10/NET4536 0 0.176433f
c_330 XI10/NET4752 0 0.176433f
c_331 XI10/NET4460 0 0.176433f
c_332 XI10/NET4700 0 0.176433f
c_333 XI10/NET5416 0 0.176433f
c_334 XI10/NET5200 0 0.176433f
c_335 XI10/NET4292 0 0.176433f
c_336 XI10/NET5176 0 0.176433f
c_337 XI10/NET2100 0 0.176433f
c_338 XI10/NET2316 0 0.176433f
c_339 XI10/NET2024 0 0.176433f
c_340 XI10/NET2264 0 0.176433f
c_341 XI10/NET2804 0 0.176433f
c_342 XI10/NET02612 0 0.176433f
c_343 XI10/NET2880 0 0.176433f
c_344 XI10/NET2548 0 0.176433f
c_345 XI10/NET5596 0 0.176433f
c_346 XI10/NET1836 0 0.176433f
c_347 XI10/NET5520 0 0.176433f
c_348 XI10/NET1796 0 0.176433f
c_349 XI10/NET3052 0 0.176433f
c_350 XI10/NET3268 0 0.176433f
c_351 XI10/NET1952 0 0.176433f
c_352 XI10/NET3216 0 0.176433f
c_353 XI10/NET3680 0 0.18051f
c_354 XI10/NET3632 0 0.176433f
c_355 XI10/NET3888 0 0.176433f
c_356 XI10/NET4908 0 0.176433f
c_357 XI10/NET4136 0 0.176433f
c_358 XI10/NET4204 0 0.176433f
c_359 XI10/NET3928 0 0.176433f
c_360 XI10/NET3552 0 0.176433f
c_361 XI10/NET4604 0 0.18066f
c_362 XI10/NET4672 0 0.176433f
c_363 XI10/NET4412 0 0.176433f
c_364 XI10/NET4828 0 0.176433f
c_365 XI10/NET5348 0 0.176433f
c_366 XI10/NET5268 0 0.176433f
c_367 XI10/NET4356 0 0.176433f
c_368 XI10/NET5124 0 0.176433f
c_369 XI10/NET2168 0 0.18066f
c_370 XI10/NET2236 0 0.176433f
c_371 XI10/NET2440 0 0.176433f
c_372 XI10/NET2392 0 0.176433f
c_373 XI10/NET2736 0 0.176433f
c_374 XI10/NET2656 0 0.176433f
c_375 XI10/NET2924 0 0.176433f
c_376 XI10/NET2512 0 0.176433f
c_377 XI10/NET5664 0 0.18066f
c_378 XI10/NET5736 0 0.176433f
c_379 XI10/NET3320 0 0.176433f
c_380 XI10/NET1760 0 0.176433f
c_381 XI10/NET3120 0 0.176433f
c_382 XI10/NET3188 0 0.176433f
c_383 XI10/NET1904 0 0.176433f
c_384 XI10/NET3384 0 0.176433f
c_385 XI10/NET3736 0 0.176433f
c_386 XI10/NET5012 0 0.176433f
c_387 XI10/NET3812 0 0.176433f
c_388 XI10/NET3792 0 0.176433f
c_389 XI10/NET4056 0 0.176433f
c_390 XI10/NET3448 0 0.176433f
c_391 XI10/NET3980 0 0.176433f
c_392 XI10/NET3516 0 0.176433f
c_393 XI10/NET4524 0 0.176433f
c_394 XI10/NET4740 0 0.176433f
c_395 XI10/NET4448 0 0.176433f
c_396 XI10/NET4660 0 0.176433f
c_397 XI10/NET5404 0 0.176433f
c_398 XI10/NET5188 0 0.176433f
c_399 XI10/NET4280 0 0.176433f
c_400 XI10/NET5164 0 0.176433f
c_401 XI10/NET2088 0 0.176433f
c_402 XI10/NET2304 0 0.176433f
c_403 XI10/NET2012 0 0.176433f
c_404 XI10/NET2224 0 0.176433f
c_405 XI10/NET2792 0 0.176433f
c_406 XI10/NET02600 0 0.176433f
c_407 XI10/NET2868 0 0.176433f
c_408 XI10/NET2480 0 0.176433f
c_409 XI10/NET5584 0 0.176433f
c_410 XI10/NET1824 0 0.176433f
c_411 XI10/NET5508 0 0.176433f
c_412 XI10/NET1728 0 0.176433f
c_413 XI10/NET3040 0 0.176433f
c_414 XI10/NET3256 0 0.176433f
c_415 XI10/NET1940 0 0.176433f
c_416 XI10/NET3176 0 0.176433f
c_417 XI10/NET3668 0 0.18051f
c_418 XI10/NET3624 0 0.176433f
c_419 XI10/NET3876 0 0.176433f
c_420 XI10/NET3800 0 0.176433f
c_421 XI10/NET4124 0 0.176433f
c_422 XI10/NET4188 0 0.176433f
c_423 XI10/NET3584 0 0.176433f
c_424 XI10/NET3540 0 0.176433f
c_425 XI10/NET4592 0 0.18066f
c_426 XI10/NET4656 0 0.176433f
c_427 XI10/NET4400 0 0.176433f
c_428 XI10/NET4580 0 0.176433f
c_429 XI10/NET5336 0 0.176433f
c_430 XI10/NET5256 0 0.176433f
c_431 XI10/NET4344 0 0.176433f
c_432 XI10/NET5108 0 0.176433f
c_433 XI10/NET2156 0 0.18066f
c_434 XI10/NET2220 0 0.176433f
c_435 XI10/NET2424 0 0.176433f
c_436 XI10/NET2144 0 0.176433f
c_437 XI10/NET2724 0 0.176433f
c_438 XI10/NET2644 0 0.176433f
c_439 XI10/NET2500 0 0.176433f
c_440 XI10/NET2496 0 0.176433f
c_441 XI10/NET5652 0 0.18066f
c_442 XI10/NET5720 0 0.176433f
c_443 XI10/NET1748 0 0.176433f
c_444 XI10/NET1744 0 0.176433f
c_445 XI10/NET3108 0 0.176433f
c_446 XI10/NET3172 0 0.176433f
c_447 XI10/NET1892 0 0.176433f
c_448 XI10/NET3096 0 0.176433f
c_449 XI10/NET3788 0 0.176433f
c_450 XI10/NET5004 0 0.176433f
c_451 XI10/NET3804 0 0.176433f
c_452 XI10/NET3644 0 0.176433f
c_453 XI10/NET4048 0 0.176433f
c_454 XI10/NET3444 0 0.176433f
c_455 XI10/NET3976 0 0.176433f
c_456 XI10/NET3504 0 0.176433f
c_457 XI10/NET4516 0 0.176433f
c_458 XI10/NET4736 0 0.176433f
c_459 XI10/NET4444 0 0.176433f
c_460 XI10/NET4512 0 0.176433f
c_461 XI10/NET5400 0 0.176433f
c_462 XI10/NET5180 0 0.176433f
c_463 XI10/NET4272 0 0.176433f
c_464 XI10/NET5160 0 0.176433f
c_465 XI10/NET2080 0 0.176433f
c_466 XI10/NET2300 0 0.176433f
c_467 XI10/NET2008 0 0.176433f
c_468 XI10/NET2076 0 0.176433f
c_469 XI10/NET2788 0 0.176433f
c_470 XI10/NET02592 0 0.176433f
c_471 XI10/NET2860 0 0.176433f
c_472 XI10/NET2464 0 0.176433f
c_473 XI10/NET5576 0 0.176433f
c_474 XI10/NET1816 0 0.176433f
c_475 XI10/NET5504 0 0.176433f
c_476 XI10/NET1712 0 0.176433f
c_477 XI10/NET3032 0 0.176433f
c_478 XI10/NET3252 0 0.176433f
c_479 XI10/NET1936 0 0.176433f
c_480 XI10/NET3028 0 0.176433f
c_481 XI10/NET3664 0 0.140391f
c_482 XI10/NET3608 0 0.136314f
c_483 XI10/NET3868 0 0.136314f
c_484 XI10/NET3724 0 0.136314f
c_485 XI10/NET4116 0 0.136314f
c_486 XI10/NET4184 0 0.136314f
c_487 XI10/NET3568 0 0.136314f
c_488 XI10/NET3536 0 0.136314f
c_489 XI10/NET4584 0 0.138908f
c_490 XI10/NET4652 0 0.136314f
c_491 XI10/NET4396 0 0.136314f
c_492 XI10/NET4504 0 0.136314f
c_493 XI10/NET5332 0 0.136314f
c_494 XI10/NET5244 0 0.136314f
c_495 XI10/NET4336 0 0.136314f
c_496 XI10/NET4268 0 0.136314f
c_497 XI10/NET2148 0 0.138908f
c_498 XI10/NET2216 0 0.136314f
c_499 XI10/NET2000 0 0.136314f
c_500 XI10/NET2068 0 0.136314f
c_501 XI10/NET2720 0 0.136314f
c_502 XI10/NET2632 0 0.136314f
c_503 XI10/NET2484 0 0.136314f
c_504 XI10/NET2472 0 0.136314f
c_505 XI10/NET5644 0 0.138908f
c_506 XI10/NET5716 0 0.136314f
c_507 XI10/NET1732 0 0.136314f
c_508 XI10/NET1720 0 0.136314f
c_509 XI10/NET3100 0 0.136314f
c_510 XI10/NET3168 0 0.136314f
c_511 XI10/NET1888 0 0.136314f
c_512 XI10/NET1996 0 0.136314f
*
.include "Final_all_v1.pex.spi.FINAL_ALL_V1.pxi"
*
.ends
*
*
