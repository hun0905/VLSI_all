* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT mos_unit
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nor_small 1 2 3 4 5 7 8
** N=8 EP=7 IP=12 FDC=4
M0 2 1 5 2 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-1665 $Y=1620 $D=0
M1 5 3 2 2 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-205 $Y=1620 $D=0
M2 6 3 4 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-5290 $Y=1620 $D=1
M3 5 1 6 8 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-3830 $Y=1620 $D=1
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=8
X0 1 2 3 6 7 9 10 nor_small $T=0 0 0 0 $X=-22995 $Y=1285
X1 4 2 5 6 8 11 12 nor_small $T=0 1525 0 0 $X=-22995 $Y=2810
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21
** N=21 EP=21 IP=24 FDC=16
X0 1 3 4 2 5 9 10 11 14 15 16 17 ICV_1 $T=0 0 0 0 $X=-22995 $Y=1285
X1 6 3 5 7 8 9 12 13 18 19 20 21 ICV_1 $T=0 3050 0 0 $X=-22995 $Y=4335
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38
** N=38 EP=38 IP=42 FDC=32
X0 1 2 5 6 7 3 4 8 14 15 16 17 18 23 24 25 26 27 28 29
+ 30
+ ICV_2 $T=0 0 0 0 $X=-22995 $Y=1285
X1 9 10 5 8 8 11 12 13 14 19 20 21 22 31 32 33 34 35 36 37
+ 38
+ ICV_2 $T=0 6100 0 0 $X=-22995 $Y=7385
.ENDS
***************************************
.SUBCKT inv_small 1 2 3 4 5 6 7
** N=7 EP=7 IP=12 FDC=4
M0 4 2 1 4 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=1485 $Y=-590 $D=0
M1 1 2 3 5 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-2060 $Y=-590 $D=1
M2 3 2 1 6 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-1370 $Y=-590 $D=1
M3 1 2 3 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-680 $Y=-590 $D=1
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=8
X0 2 1 5 6 7 8 9 inv_small $T=0 0 0 0 $X=-3295 $Y=-1110
X1 4 3 5 6 10 11 12 inv_small $T=0 1960 0 0 $X=-3295 $Y=850
.ENDS
***************************************
.SUBCKT nand_small_hw4 1 2 3 4 5 6 9 10 11 12 13 14 15 16 17
** N=17 EP=15 IP=36 FDC=12
M0 7 2 3 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=3610 $Y=-1710 $D=0
M1 8 4 7 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=5105 $Y=-1710 $D=0
M2 5 1 8 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=6565 $Y=-1710 $D=0
M3 3 1 6 9 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-5610 $Y=-1710 $D=1
M4 6 1 3 10 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-4920 $Y=-1710 $D=1
M5 3 1 6 11 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-4230 $Y=-1710 $D=1
M6 3 4 6 12 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-2770 $Y=-1710 $D=1
M7 6 4 3 13 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-2080 $Y=-1710 $D=1
M8 3 4 6 14 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=-1390 $Y=-1710 $D=1
M9 3 2 6 15 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=70 $Y=-1710 $D=1
M10 6 2 3 16 P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=760 $Y=-1710 $D=1
M11 3 2 6 17 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=1450 $Y=-1710 $D=1
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26
** N=26 EP=26 IP=30 FDC=24
X0 3 1 7 2 4 6 9 10 11 12 13 14 15 16 17 nand_small_hw4 $T=0 0 0 0 $X=-22630 $Y=-2570
X1 5 1 8 2 4 6 18 19 20 21 22 23 24 25 26 nand_small_hw4 $T=0 3440 0 0 $X=-22630 $Y=870
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47
** N=47 EP=47 IP=52 FDC=48
X0 1 2 3 5 4 7 8 9 12 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29
+ ICV_5 $T=0 0 0 0 $X=-22630 $Y=-2570
X1 1 6 3 5 4 7 10 11 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47
+ ICV_5 $T=0 6880 0 0 $X=-22630 $Y=4310
.ENDS
***************************************
.SUBCKT hw4_decoder in<5> in<4> in<3> in<2> in<1> in<0> VDD VSS OUT<55> OUT<0> OUT<34> OUT<33> OUT<12> OUT<11> OUT<2> OUT<1> OUT<38> OUT<37> OUT<36> OUT<35>
+ OUT<16> OUT<15> OUT<14> OUT<13> OUT<63> OUT<62> OUT<61> OUT<60> OUT<59> OUT<58> OUT<57> OUT<56> OUT<54> OUT<53> OUT<52> OUT<51> OUT<50> OUT<49> OUT<48> OUT<47>
+ OUT<46> OUT<45> OUT<44> OUT<43> OUT<42> OUT<41> OUT<40> OUT<39> OUT<32> OUT<31> OUT<30> OUT<29> OUT<28> OUT<27> OUT<26> OUT<25> OUT<24> OUT<23> OUT<22> OUT<21>
+ OUT<20> OUT<19> OUT<18> OUT<17> OUT<10> OUT<9> OUT<8> OUT<7> OUT<6> OUT<5> OUT<4> OUT<3>
** N=94 EP=72 IP=546 FDC=472
X0 20 VSS 28 VDD OUT<55> VDD VDD nor_small $T=22910 101150 0 0 $X=-85 $Y=102435
X1 18 VSS 13 VDD OUT<0> VDD VDD nor_small $T=22910 187670 0 0 $X=-85 $Y=188955
X2 16 VSS 27 19 27 VDD OUT<34> OUT<33> VDD VDD VDD VDD ICV_1 $T=22910 134080 0 0 $X=-85 $Y=135365
X3 22 VSS 15 14 15 VDD OUT<12> OUT<11> VDD VDD VDD VDD ICV_1 $T=22910 168500 0 0 $X=-85 $Y=169785
X4 16 VSS 13 19 13 VDD OUT<2> OUT<1> VDD VDD VDD VDD ICV_1 $T=22910 184620 0 0 $X=-85 $Y=185905
X5 21 17 VSS 27 27 22 14 27 VDD OUT<38> OUT<37> OUT<36> OUT<35> VDD VDD VDD VDD VDD VDD VDD
+ VDD
+ ICV_2 $T=22910 127980 0 0 $X=-85 $Y=129265
X6 18 20 VSS 24 15 21 17 15 VDD OUT<16> OUT<15> OUT<14> OUT<13> VDD VDD VDD VDD VDD VDD VDD
+ VDD
+ ICV_2 $T=22910 162400 0 0 $X=-85 $Y=163685
X7 20 21 17 22 VSS 23 23 23 14 16 19 18 23 VDD OUT<63> OUT<62> OUT<61> OUT<60> OUT<59> OUT<58>
+ OUT<57> OUT<56> VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ ICV_3 $T=22910 88950 0 0 $X=-85 $Y=90235
X8 21 17 22 14 VSS 28 28 28 16 19 18 20 25 VDD OUT<54> OUT<53> OUT<52> OUT<51> OUT<50> OUT<49>
+ OUT<48> OUT<47> VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ ICV_3 $T=22910 103580 0 0 $X=-85 $Y=104865
X9 21 17 22 14 VSS 25 25 25 16 19 18 20 27 VDD OUT<46> OUT<45> OUT<44> OUT<43> OUT<42> OUT<41>
+ OUT<40> OUT<39> VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ ICV_3 $T=22910 115780 0 0 $X=-85 $Y=117065
X10 18 20 21 17 VSS 27 26 26 22 14 16 19 26 VDD OUT<32> OUT<31> OUT<30> OUT<29> OUT<28> OUT<27>
+ OUT<26> OUT<25> VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ ICV_3 $T=22910 138000 0 0 $X=-85 $Y=139285
X11 18 20 21 17 VSS 26 24 24 22 14 16 19 24 VDD OUT<24> OUT<23> OUT<22> OUT<21> OUT<20> OUT<19>
+ OUT<18> OUT<17> VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ ICV_3 $T=22910 150200 0 0 $X=-85 $Y=151485
X12 16 19 18 20 VSS 15 15 13 21 17 22 14 13 VDD OUT<10> OUT<9> OUT<8> OUT<7> OUT<6> OUT<5>
+ OUT<4> OUT<3> VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ ICV_3 $T=22910 172420 0 0 $X=-85 $Y=173705
X13 6 in<3> VDD VSS VDD VDD VDD inv_small $T=-41095 184355 0 0 $X=-44390 $Y=183245
X14 12 in<0> VDD VSS VDD VDD VDD inv_small $T=-20335 184355 0 0 $X=-23630 $Y=183245
X15 in<5> 4 in<4> 5 VDD VSS VDD VDD VDD VDD VDD VDD ICV_4 $T=-41095 180435 0 0 $X=-44390 $Y=179325
X16 in<2> 10 in<1> 11 VDD VSS VDD VDD VDD VDD VDD VDD ICV_4 $T=-20335 180435 0 0 $X=-23630 $Y=179325
X17 in<2> in<1> in<0> 12 VSS 11 VDD 20 21 17 22 VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD
+ ICV_6 $T=-19595 137695 0 0 $X=-42225 $Y=135125
X18 10 in<1> in<0> 12 VSS 11 VDD 14 16 19 18 VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD
+ ICV_6 $T=-19595 152325 0 0 $X=-42225 $Y=149755
X19 in<5> in<4> in<3> 6 VSS 5 VDD 23 28 25 27 VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD
+ ICV_6 $T=-19525 109305 0 0 $X=-42155 $Y=106735
X20 4 in<4> in<3> 6 VSS 5 VDD 26 24 15 13 VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD VDD VDD VDD VDD
+ ICV_6 $T=-19525 123935 0 0 $X=-42155 $Y=121365
.ENDS
***************************************
