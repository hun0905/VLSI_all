* File: hw3_part2.pex.spi
* Created: Sat Nov 27 18:15:55 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw3_part2.pex.spi.pex"
.subckt hw3_part2  VSS C NET14 VDD !C D Q !Q
* 
* !Q	!Q
* Q	Q
* D	D
* !C	!C
* VDD	VDD
* NET14	NET14
* C	C
* VSS	VSS
MM0 N_NET18_MM0_d N_C_MM0_g N_NET13_MM0_s N_VDD_XI0/MM6_b P_18 L=1.8e-07
+ W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
MM3 N_NET5_MM3_d N_!C_MM3_g N_NET14_MM3_s N_VDD_MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
MM2 N_NET18_MM2_d N_!C_MM2_g N_NET13_MM2_s N_VSS_MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM1 N_NET5_MM1_d N_C_MM1_g N_NET14_MM1_s N_VSS_MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0/MM6 N_NET18_XI0/MM6_d N_D_XI0/MM6_g N_VDD_XI0/MM6_s N_VDD_XI0/MM6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0/MM10 N_NET18_XI0/MM10_d N_D_XI0/MM10_g N_VSS_XI0/MM10_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1/MM6 N_NET14_XI1/MM6_d N_NET13_XI1/MM6_g N_VDD_XI1/MM6_s N_VDD_XI0/MM6_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1/MM10 N_NET14_XI1/MM10_d N_NET13_XI1/MM10_g N_VSS_XI1/MM10_s N_VSS_MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI4/MM6 N_Q_XI4/MM6_d N_NET1_XI4/MM6_g N_VDD_XI4/MM6_s N_VDD_XI4/MM6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI4/MM10 N_Q_XI4/MM10_d N_NET1_XI4/MM10_g N_VSS_XI4/MM10_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI3/MM6 N_NET1_XI3/MM6_d N_NET5_XI3/MM6_g N_VDD_XI3/MM6_s N_VDD_XI3/MM6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI3/MM10 N_NET1_XI3/MM10_d N_NET5_XI3/MM10_g N_VSS_XI3/MM10_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI2/MM6 N_!Q_XI2/MM6_d N_NET5_XI2/MM6_g N_VDD_XI2/MM6_s N_VDD_XI2/MM6_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI2/MM10 N_!Q_XI2/MM10_d N_NET5_XI2/MM10_g N_VSS_XI2/MM10_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/MM1 N_NET13_XI5/MM1_d N_NET14_XI5/MM1_g N_XI5/NET12_XI5/MM1_s
+ N_VDD_XI5/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI5/MM0 N_XI5/NET12_XI5/MM0_d N_!C_XI5/MM0_g N_VDD_XI5/MM0_s N_VDD_XI5/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI5/MM2 N_NET13_XI5/MM2_d N_NET14_XI5/MM2_g N_XI5/NET5_XI5/MM2_s N_VSS_MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/MM3 N_XI5/NET5_XI5/MM3_d N_C_XI5/MM3_g N_VSS_XI5/MM3_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI6/MM1 N_NET5_XI6/MM1_d N_NET1_XI6/MM1_g N_XI6/NET12_XI6/MM1_s N_VDD_XI6/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI6/MM0 N_XI6/NET12_XI6/MM0_d N_C_XI6/MM0_g N_VDD_XI6/MM0_s N_VDD_XI6/MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI6/MM2 N_NET5_XI6/MM2_d N_NET1_XI6/MM2_g N_XI6/NET5_XI6/MM2_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI6/MM3 N_XI6/NET5_XI6/MM3_d N_!C_XI6/MM3_g N_VSS_XI6/MM3_s N_VSS_MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
*
.include "hw3_part2.pex.spi.HW3_PART2.pxi"
*
.ends
*
*
