* File: hw2_part2_1.pex.spi
* Created: Fri Nov 12 00:28:27 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw2_part2_1.pex.spi.pex"
.subckt hw2_part2_1  IN OUT OUT2 OUT3 OUT4 VSS VDD OUT5
* 
* OUT5	OUT5
* VDD	VDD
* VSS	VSS
* OUT4	OUT4
* OUT3	OUT3
* OUT2	OUT2
* OUT	OUT
* IN	IN
MM8 N_OUT3_MM8_d N_OUT2_MM8_g N_VSS_MM8_s N_VSS_MM10_b N_18 L=1.8e-07 W=2.5e-06
+ AD=1.225e-12 AS=1.225e-12 PD=3.48e-06 PS=3.48e-06
MM9 N_OUT4_MM9_d N_OUT3_MM9_g N_VSS_MM9_s N_VSS_MM10_b N_18 L=1.8e-07 W=2.5e-06
+ AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM9@5 N_OUT4_MM9@5_d N_OUT3_MM9@5_g N_VSS_MM9@5_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM9@4 N_OUT4_MM9@4_d N_OUT3_MM9@4_g N_VSS_MM9@4_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM9@3 N_OUT4_MM9@3_d N_OUT3_MM9@3_g N_VSS_MM9@3_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM9@2 N_OUT4_MM9@2_d N_OUT3_MM9@2_g N_VSS_MM9@2_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM11 N_OUT5_MM11_d N_OUT4_MM11_g N_VSS_MM11_s N_VSS_MM10_b N_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM11@25 N_OUT5_MM11@25_d N_OUT4_MM11@25_g N_VSS_MM11@25_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@24 N_OUT5_MM11@24_d N_OUT4_MM11@24_g N_VSS_MM11@24_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@23 N_OUT5_MM11@23_d N_OUT4_MM11@23_g N_VSS_MM11@23_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@22 N_OUT5_MM11@22_d N_OUT4_MM11@22_g N_VSS_MM11@22_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@21 N_OUT5_MM11@21_d N_OUT4_MM11@21_g N_VSS_MM11@21_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@20 N_OUT5_MM11@20_d N_OUT4_MM11@20_g N_VSS_MM11@20_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@19 N_OUT5_MM11@19_d N_OUT4_MM11@19_g N_VSS_MM11@19_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@18 N_OUT5_MM11@18_d N_OUT4_MM11@18_g N_VSS_MM11@18_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@17 N_OUT5_MM11@17_d N_OUT4_MM11@17_g N_VSS_MM11@17_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@16 N_OUT5_MM11@16_d N_OUT4_MM11@16_g N_VSS_MM11@16_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@15 N_OUT5_MM11@15_d N_OUT4_MM11@15_g N_VSS_MM11@15_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@14 N_OUT5_MM11@14_d N_OUT4_MM11@14_g N_VSS_MM11@14_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@13 N_OUT5_MM11@13_d N_OUT4_MM11@13_g N_VSS_MM11@13_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@12 N_OUT5_MM11@12_d N_OUT4_MM11@12_g N_VSS_MM11@12_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@11 N_OUT5_MM11@11_d N_OUT4_MM11@11_g N_VSS_MM11@11_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@10 N_OUT5_MM11@10_d N_OUT4_MM11@10_g N_VSS_MM11@10_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@9 N_OUT5_MM11@9_d N_OUT4_MM11@9_g N_VSS_MM11@9_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@8 N_OUT5_MM11@8_d N_OUT4_MM11@8_g N_VSS_MM11@8_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@7 N_OUT5_MM11@7_d N_OUT4_MM11@7_g N_VSS_MM11@7_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@6 N_OUT5_MM11@6_d N_OUT4_MM11@6_g N_VSS_MM11@6_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@5 N_OUT5_MM11@5_d N_OUT4_MM11@5_g N_VSS_MM11@5_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@4 N_OUT5_MM11@4_d N_OUT4_MM11@4_g N_VSS_MM11@4_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@3 N_OUT5_MM11@3_d N_OUT4_MM11@3_g N_VSS_MM11@3_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM11@2 N_OUT5_MM11@2_d N_OUT4_MM11@2_g N_VSS_MM11@2_s N_VSS_MM10_b N_18
+ L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM10 N_OUT_MM10_d N_IN_MM10_g N_VSS_MM10_s N_VSS_MM10_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM4 N_OUT2_MM4_d N_OUT_MM4_g N_VSS_MM4_s N_VSS_MM10_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM7 N_OUT5_MM7_d N_OUT4_MM7_g N_VDD_MM7_s N_VDD_MM6_b P_18 L=1.8e-07 W=2.5e-06
+ AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06
MM7@25 N_OUT5_MM7@25_d N_OUT4_MM7@25_g N_VDD_MM7@25_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@24 N_OUT5_MM7@24_d N_OUT4_MM7@24_g N_VDD_MM7@24_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@23 N_OUT5_MM7@23_d N_OUT4_MM7@23_g N_VDD_MM7@23_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@22 N_OUT5_MM7@22_d N_OUT4_MM7@22_g N_VDD_MM7@22_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@21 N_OUT5_MM7@21_d N_OUT4_MM7@21_g N_VDD_MM7@21_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@20 N_OUT5_MM7@20_d N_OUT4_MM7@20_g N_VDD_MM7@20_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@19 N_OUT5_MM7@19_d N_OUT4_MM7@19_g N_VDD_MM7@19_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@18 N_OUT5_MM7@18_d N_OUT4_MM7@18_g N_VDD_MM7@18_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@17 N_OUT5_MM7@17_d N_OUT4_MM7@17_g N_VDD_MM7@17_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@16 N_OUT5_MM7@16_d N_OUT4_MM7@16_g N_VDD_MM7@16_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@15 N_OUT5_MM7@15_d N_OUT4_MM7@15_g N_VDD_MM7@15_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@14 N_OUT5_MM7@14_d N_OUT4_MM7@14_g N_VDD_MM7@14_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@13 N_OUT5_MM7@13_d N_OUT4_MM7@13_g N_VDD_MM7@13_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@12 N_OUT5_MM7@12_d N_OUT4_MM7@12_g N_VDD_MM7@12_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@11 N_OUT5_MM7@11_d N_OUT4_MM7@11_g N_VDD_MM7@11_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@10 N_OUT5_MM7@10_d N_OUT4_MM7@10_g N_VDD_MM7@10_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@9 N_OUT5_MM7@9_d N_OUT4_MM7@9_g N_VDD_MM7@9_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@8 N_OUT5_MM7@8_d N_OUT4_MM7@8_g N_VDD_MM7@8_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@7 N_OUT5_MM7@7_d N_OUT4_MM7@7_g N_VDD_MM7@7_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@6 N_OUT5_MM7@6_d N_OUT4_MM7@6_g N_VDD_MM7@6_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@5 N_OUT5_MM7@5_d N_OUT4_MM7@5_g N_VDD_MM7@5_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@4 N_OUT5_MM7@4_d N_OUT4_MM7@4_g N_VDD_MM7@4_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@3 N_OUT5_MM7@3_d N_OUT4_MM7@3_g N_VDD_MM7@3_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07
MM7@2 N_OUT5_MM7@2_d N_OUT4_MM7@2_g N_VDD_MM7@2_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07
MM6 N_OUT_MM6_d N_IN_MM6_g N_VDD_MM6_s N_VDD_MM6_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM0 N_OUT2_MM0_d N_OUT_MM0_g N_VDD_MM0_s N_VDD_MM6_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM3 N_OUT3_MM3_d N_OUT2_MM3_g N_VDD_MM3_s N_VDD_MM6_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
MM5 N_OUT4_MM5_d N_OUT3_MM5_g N_VDD_MM5_s N_VDD_MM6_b P_18 L=1.8e-07 W=1.85e-06
+ AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
MM5@5 N_OUT4_MM5@5_d N_OUT3_MM5@5_g N_VDD_MM5@5_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM5@4 N_OUT4_MM5@4_d N_OUT3_MM5@4_g N_VDD_MM5@4_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM5@3 N_OUT4_MM5@3_d N_OUT3_MM5@3_g N_VDD_MM5@3_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=1.85e-06 AD=4.7175e-13 AS=4.7175e-13 PD=5.1e-07 PS=5.1e-07
MM5@2 N_OUT4_MM5@2_d N_OUT3_MM5@2_g N_VDD_MM5@2_s N_VDD_MM6_b P_18 L=1.8e-07
+ W=1.85e-06 AD=9.065e-13 AS=4.7175e-13 PD=2.83e-06 PS=5.1e-07
*
.include "hw2_part2_1.pex.spi.HW2_PART2_1.pxi"
*
.ends
*
*
