* File: hw5_SA.pex.spi
* Created: Tue Dec 28 00:50:29 2021
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "hw5_SA.pex.spi.pex"
.subckt hw5  SON SO COM VSS INN EN VDD INP
.PARAM VTH = AGAUSS(0,0.072,6) 
* INP	INP
* VDD	VDD
* EN	EN
* INN	INN
* VSS	VSS
* COM	COM
* SO	SO
* SON	SON
MM16 N_NET093_MM16_d N_INN_MM16_g N_COM_MM16_s N_VSS_MM16_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM15 N_SO_MM15_d N_SON_MM15_g N_NET093_MM15_s N_VSS_MM16_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM19 N_COM_MM19_d N_EN_MM19_g N_VSS_MM19_s N_VSS_MM16_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 delvto=VTH
MM19@3 N_COM_MM19@3_d N_EN_MM19@3_g N_VSS_MM19@3_s N_VSS_MM16_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 delvto=VTH
MM19@2 N_COM_MM19@2_d N_EN_MM19@2_g N_VSS_MM19@2_s N_VSS_MM16_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 delvto=VTH
MM17 N_SON_MM17_d N_SO_MM17_g N_NET089_MM17_s N_VSS_MM16_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM18 N_NET089_MM18_d N_INP_MM18_g N_COM_MM18_s N_VSS_MM16_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM12 N_SO_MM12_d N_SON_MM12_g N_VDD_MM12_s N_VDD_MM12_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM11 N_SO_MM11_d N_EN_MM11_g N_VDD_MM11_s N_VDD_MM12_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM9 N_SON_MM9_d N_EN_MM9_g N_VDD_MM9_s N_VDD_MM12_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
MM13 N_SON_MM13_d N_SO_MM13_g N_VDD_MM13_s N_VDD_MM12_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 delvto=VTH
*
.include "hw5_SA.pex.spi.HW5_SA.pxi"
*
.ends
*
*
