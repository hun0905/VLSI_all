************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: nand3
* View Name:     schematic
* Netlisted on:  Oct 30 21:11:47 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    nand3
* View Name:    schematic
************************************************************************

.SUBCKT nand3 A B C OUT VDD VSS
*.PININFO A:I B:I C:I OUT:O VDD:B VSS:B
MM6 net6 C VSS VSS NM W=8u L=180.00n m=1
MM5 net10 B net6 VSS NM W=8u L=180.00n m=1
MM4 OUT A net10 VSS NM W=8u L=180.00n m=1
MM2 OUT C VDD VDD PM W=1.65u L=180.00n m=1
MM1 OUT A VDD VDD PM W=13.2u L=180.00n m=1
MM0 OUT B VDD VDD PM W=1.65u L=180.00n m=1
.ENDS

