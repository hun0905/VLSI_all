************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: hw2_part2_1
* View Name:     schematic
* Netlisted on:  Nov 11 15:36:17 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    hw2_part2_1
* View Name:    schematic
************************************************************************

.SUBCKT hw2_part2_1 IN OUT OUT2 OUT3 OUT4 OUT5 VDD VSS
*.PININFO IN:I OUT5:O OUT:B OUT2:B OUT3:B OUT4:B VDD:B VSS:B
MM11 OUT5 OUT4 VSS VSS NM W=2.5u L=180.00n m=20
MM8 OUT3 OUT2 VSS VSS NM W=500.0n L=180.00n m=1
MM9 OUT4 OUT3 VSS VSS NM W=500.0n L=180.00n m=5
MM10 OUT IN VSS VSS NM W=500.0n L=180.00n m=1
MM4 OUT2 OUT VSS VSS NM W=500.0n L=180.00n m=1
MM7 OUT5 OUT4 VDD VDD PM W=2.5u L=180.00n m=25
MM3 OUT3 OUT2 VDD VDD PM W=1.85u L=180.00n m=1
MM5 OUT4 OUT3 VDD VDD PM W=1.85u L=180.00n m=5
MM6 OUT IN VDD VDD PM W=1.85u L=180.00n m=1
MM0 OUT2 OUT VDD VDD PM W=1.85u L=180.00n m=1
.ENDS

