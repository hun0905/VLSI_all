************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: YMUX
* View Name:     schematic
* Netlisted on:  Jan 12 01:21:35 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter IN OUT VDD VSS
*.PININFO IN:I OUT:B VDD:B VSS:B
MM10 OUT IN VSS VSS N_18 W=500.0n L=180.00n m=1
MM6 OUT IN VDD VDD P_18 W=2u L=180.00n m=1
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG BL OUT SEL VDD VSS
*.PININFO BL:I SEL:I VDD:I VSS:I OUT:O
XI1 SEL net40 VDD VSS / inverter
MM1 BL SEL OUT VSS N_18 W=500.0n L=180.00n
MM0 BL net40 OUT VDD P_18 W=1.5u L=180.00n
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    YMUX
* View Name:    schematic
************************************************************************

.SUBCKT YMUX BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> Dout VDD VSS 
+ Ysel<0> Ysel<1> Ysel<2> Ysel<3> Ysel<4> Ysel<5> Ysel<6> Ysel<7>
*.PININFO BL<0>:I BL<1>:I BL<2>:I BL<3>:I BL<4>:I BL<5>:I BL<6>:I BL<7>:I 
*.PININFO Ysel<0>:I Ysel<1>:I Ysel<2>:I Ysel<3>:I Ysel<4>:I Ysel<5>:I 
*.PININFO Ysel<6>:I Ysel<7>:I Dout:O VDD:B VSS:B
XI15 BL<4> Dout Ysel<4> VDD VSS / TG
XI18 BL<7> Dout Ysel<7> VDD VSS / TG
XI19 BL<3> Dout Ysel<3> VDD VSS / TG
XI20 BL<2> Dout Ysel<2> VDD VSS / TG
XI21 BL<1> Dout Ysel<1> VDD VSS / TG
XI22 BL<0> Dout Ysel<0> VDD VSS / TG
XI16 BL<5> Dout Ysel<5> VDD VSS / TG
XI17 BL<6> Dout Ysel<6> VDD VSS / TG
.ENDS

