* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT mos_unit2
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT mos_unit
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Final_SA 1 2 3 4 5 6 7
** N=10 EP=7 IP=40 FDC=12
M0 9 4 8 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-2175 $Y=-410 $D=0
M1 5 3 8 5 N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=-1310 $Y=-1590 $D=0
M2 2 1 9 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-715 $Y=-410 $D=0
M3 8 3 5 5 N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=-620 $Y=-1590 $D=0
M4 5 3 8 5 N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=70 $Y=-1590 $D=0
M5 10 2 1 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=745 $Y=-410 $D=0
M6 8 3 5 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=760 $Y=-1590 $D=0
M7 8 6 10 5 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=2205 $Y=-410 $D=0
M8 2 3 7 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-2175 $Y=1410 $D=1
M9 2 1 7 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-715 $Y=1410 $D=1
M10 7 2 1 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=745 $Y=1410 $D=1
M11 7 3 1 7 P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=2205 $Y=1410 $D=1
.ENDS
***************************************
.SUBCKT final_mos_unit
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT inv_final 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 2 2 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-65 $Y=-2195 $D=0
M1 4 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-65 $Y=-490 $D=1
.ENDS
***************************************
.SUBCKT final_and 1 2 3 4 5
** N=7 EP=5 IP=28 FDC=6
M0 7 2 4 4 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=8825 $Y=670 $D=0
M1 6 1 7 4 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=8825 $Y=2130 $D=0
M2 6 2 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10465 $Y=670 $D=1
M3 6 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10465 $Y=2130 $D=1
X12 6 4 3 5 inv_final $T=14700 2115 0 0 $X=13540 $Y=-1150
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X0 1 2 3 4 inv_final $T=0 0 0 0 $X=-1160 $Y=-3265
X1 4 2 3 5 inv_final $T=1600 0 0 0 $X=440 $Y=-3265
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5
** N=7 EP=5 IP=10 FDC=8
X0 1 2 3 6 7 ICV_1 $T=0 0 0 0 $X=-1160 $Y=-3265
X1 7 2 3 4 5 ICV_1 $T=3200 0 0 0 $X=2040 $Y=-3265
.ENDS
***************************************
.SUBCKT inv_1u5_0u5 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 2 2 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-65 $Y=-2195 $D=0
M1 4 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-65 $Y=-490 $D=1
.ENDS
***************************************
.SUBCKT ICV_3
** N=6 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT nand4_final
** N=9 EP=0 IP=24 FDC=0
.ENDS
***************************************
.SUBCKT Ydecoder_final 1 2 3 4 5 6 7 8 9 10 11 12 13
** N=40 EP=13 IP=84 FDC=70
M0 17 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=-1665 $D=0
M1 21 3 17 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=-205 $D=0
M2 25 2 21 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=1255 $D=0
M3 4 14 25 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=2715 $D=0
M4 18 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=4355 $D=0
M5 22 16 18 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=5815 $D=0
M6 26 2 22 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=7275 $D=0
M7 5 14 26 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=8735 $D=0
M8 19 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=10375 $D=0
M9 23 3 19 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=11835 $D=0
M10 27 15 23 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=13295 $D=0
M11 6 14 27 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=14755 $D=0
M12 20 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=16395 $D=0
M13 24 16 20 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=17855 $D=0
M14 28 15 24 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=19315 $D=0
M15 7 14 28 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=9215 $Y=20775 $D=0
M16 29 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=-1645 $D=0
M17 33 3 29 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=-185 $D=0
M18 37 2 33 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=1275 $D=0
M19 8 1 37 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=2735 $D=0
M20 30 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=4375 $D=0
M21 34 16 30 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=5835 $D=0
M22 38 2 34 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=7295 $D=0
M23 9 1 38 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=8755 $D=0
M24 31 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=10395 $D=0
M25 35 3 31 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=11855 $D=0
M26 39 15 35 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=13315 $D=0
M27 10 1 39 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=14775 $D=0
M28 32 12 13 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=16415 $D=0
M29 36 16 32 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=17875 $D=0
M30 40 15 36 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=19335 $D=0
M31 11 1 40 13 N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=22140 $Y=20795 $D=0
M32 4 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=-1665 $D=1
M33 4 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=-205 $D=1
M34 4 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=1255 $D=1
M35 4 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=2715 $D=1
M36 5 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=4355 $D=1
M37 5 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=5815 $D=1
M38 5 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=7275 $D=1
M39 5 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=8735 $D=1
M40 6 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=10375 $D=1
M41 6 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=11835 $D=1
M42 6 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=13295 $D=1
M43 6 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=14755 $D=1
M44 7 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=16395 $D=1
M45 7 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=17855 $D=1
M46 7 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=19315 $D=1
M47 7 14 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=10645 $Y=20775 $D=1
M48 8 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=-1645 $D=1
M49 8 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=-185 $D=1
M50 8 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=1275 $D=1
M51 8 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=2735 $D=1
M52 9 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=4375 $D=1
M53 9 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=5835 $D=1
M54 9 2 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=7295 $D=1
M55 9 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=8755 $D=1
M56 10 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=10395 $D=1
M57 10 3 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=11855 $D=1
M58 10 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=13315 $D=1
M59 10 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=14775 $D=1
M60 11 12 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=16415 $D=1
M61 11 16 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=17875 $D=1
M62 11 15 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=19335 $D=1
M63 11 1 12 12 P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=23570 $Y=20795 $D=1
X64 3 13 12 16 inv_1u5_0u5 $T=985 1015 0 0 $X=-175 $Y=-2250
X65 2 13 12 15 inv_1u5_0u5 $T=985 7265 0 0 $X=-175 $Y=4000
X66 1 13 12 14 inv_1u5_0u5 $T=985 19305 0 0 $X=-175 $Y=16040
.ENDS
***************************************
.SUBCKT FInal_FF 1 2 3 4 5 6
** N=15 EP=6 IP=16 FDC=20
M0 9 1 7 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-2285 $Y=-2400 $D=0
M1 11 2 3 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=1670 $Y=-2400 $D=0
M2 7 12 11 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=3170 $Y=-2400 $D=0
M3 8 2 12 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=5540 $Y=-1425 $D=0
M4 13 1 3 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=9425 $Y=-2400 $D=0
M5 8 15 13 3 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10925 $Y=-2400 $D=0
M6 9 2 7 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-2285 $Y=-5120 $D=1
M7 10 1 4 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=1570 $Y=-5120 $D=1
M8 7 12 10 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=3170 $Y=-5120 $D=1
M9 8 1 12 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=5540 $Y=295 $D=1
M10 14 2 4 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=9425 $Y=-5120 $D=1
M11 8 15 14 4 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=10925 $Y=-5120 $D=1
X12 5 3 4 9 inv_1u5_0u5 $T=-2220 1570 0 0 $X=-3380 $Y=-1695
X13 7 3 4 12 inv_1u5_0u5 $T=1735 1565 0 0 $X=575 $Y=-1700
X14 8 3 4 15 inv_1u5_0u5 $T=9490 1565 0 0 $X=8330 $Y=-1700
X15 15 3 4 6 inv_1u5_0u5 $T=13725 1565 0 0 $X=12565 $Y=-1700
.ENDS
***************************************
.SUBCKT FinalProject YOUT<0> YOUT<1> YOUT<2> YOUT<3> YOUT<4> YOUT<5> YOUT<6> YOUT<7> Dout<0> SO<0> Dout<1> SO<1> VDD CLK WL_EN SAEN BL<0> BL<1> DL<0> BL<2>
+ BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> DL<1> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15> VSS X_sel<5> X_sel<2> X_sel<4> X_sel<1> X_sel<3>
+ X_sel<0> WL<63> WL<62> WL<61> WL<60> WL<59> WL<58> WL<57> WL<56> WL<55> WL<54> WL<53> WL<52> WL<51> WL<50> WL<49> WL<48> WL<47> WL<46> WL<45>
+ WL<44> WL<43> WL<42> WL<41> WL<40> WL<39> WL<38> WL<37> WL<36> WL<35> WL<34> WL<33> WL<32> WL<31> WL<30> WL<29> WL<28> WL<27> WL<26> WL<25>
+ WL<24> WL<23> WL<22> WL<21> WL<20> WL<19> WL<18> WL<17> WL<16> WL<15> WL<14> WL<13> WL<12> WL<11> WL<10> WL<9> WL<8> WL<7> WL<6> WL<5>
+ WL<4> WL<3> WL<2> WL<1> WL<0> Y_sel<0> Y_sel<2> Y_sel<1> Vref A<2> A<1> A<0> A<6> A<7> A<8> A<3> A<4> A<5>
** N=802 EP=118 IP=149 FDC=1866
M0 61 X_sel<3> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=7260 $D=0
M1 59 X_sel<4> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=19300 $D=0
M2 63 X_sel<5> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=31340 $D=0
M3 62 X_sel<0> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=55940 $D=0
M4 60 X_sel<1> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=67980 $D=0
M5 64 X_sel<2> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-66670 $Y=80020 $D=0
M6 151 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-11510 $D=0
M7 152 X_sel<3> 151 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-10050 $D=0
M8 153 X_sel<4> 152 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-8590 $D=0
M9 16 X_sel<5> 153 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-7130 $D=0
M10 154 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-5490 $D=0
M11 155 61 154 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-4030 $D=0
M12 156 X_sel<4> 155 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-2570 $D=0
M13 17 X_sel<5> 156 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=-1110 $D=0
M14 157 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=530 $D=0
M15 158 X_sel<3> 157 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=1990 $D=0
M16 159 59 158 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=3450 $D=0
M17 18 X_sel<5> 159 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=4910 $D=0
M18 160 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=6550 $D=0
M19 161 61 160 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=8010 $D=0
M20 162 59 161 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=9470 $D=0
M21 19 X_sel<5> 162 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=10930 $D=0
M22 163 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=12570 $D=0
M23 164 X_sel<3> 163 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=14030 $D=0
M24 165 X_sel<4> 164 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=15490 $D=0
M25 20 63 165 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=16950 $D=0
M26 166 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=18590 $D=0
M27 167 61 166 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=20050 $D=0
M28 168 X_sel<4> 167 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=21510 $D=0
M29 21 63 168 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=22970 $D=0
M30 169 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=24610 $D=0
M31 170 X_sel<3> 169 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=26070 $D=0
M32 171 59 170 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=27530 $D=0
M33 22 63 171 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=28990 $D=0
M34 172 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=30630 $D=0
M35 173 61 172 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=32090 $D=0
M36 174 59 173 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=33550 $D=0
M37 23 63 174 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=35010 $D=0
M38 175 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=37170 $D=0
M39 176 X_sel<0> 175 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=38630 $D=0
M40 177 X_sel<1> 176 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=40090 $D=0
M41 24 X_sel<2> 177 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=41550 $D=0
M42 178 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=43190 $D=0
M43 179 62 178 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=44650 $D=0
M44 180 X_sel<1> 179 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=46110 $D=0
M45 25 X_sel<2> 180 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=47570 $D=0
M46 181 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=49210 $D=0
M47 182 X_sel<0> 181 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=50670 $D=0
M48 183 60 182 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=52130 $D=0
M49 26 X_sel<2> 183 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=53590 $D=0
M50 184 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=55230 $D=0
M51 185 62 184 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=56690 $D=0
M52 186 60 185 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=58150 $D=0
M53 27 X_sel<2> 186 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=59610 $D=0
M54 187 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=61250 $D=0
M55 188 X_sel<0> 187 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=62710 $D=0
M56 189 X_sel<1> 188 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=64170 $D=0
M57 28 64 189 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=65630 $D=0
M58 190 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=67270 $D=0
M59 191 62 190 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=68730 $D=0
M60 192 X_sel<1> 191 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=70190 $D=0
M61 29 64 192 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=71650 $D=0
M62 193 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=73290 $D=0
M63 194 X_sel<0> 193 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=74750 $D=0
M64 195 60 194 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=76210 $D=0
M65 30 64 195 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=77670 $D=0
M66 196 WL_EN VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=79310 $D=0
M67 197 62 196 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=80770 $D=0
M68 198 60 197 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=82230 $D=0
M69 31 64 198 VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-58375 $Y=83690 $D=0
M70 WL<63> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-13505 $D=0
M71 WL<62> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-11970 $D=0
M72 WL<61> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-10435 $D=0
M73 WL<60> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-8900 $D=0
M74 WL<59> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-7365 $D=0
M75 WL<58> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-5830 $D=0
M76 WL<57> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-4295 $D=0
M77 WL<56> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-2760 $D=0
M78 WL<55> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=-1225 $D=0
M79 WL<54> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=310 $D=0
M80 WL<53> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=1845 $D=0
M81 WL<52> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=3380 $D=0
M82 WL<51> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=4915 $D=0
M83 WL<50> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=6450 $D=0
M84 WL<49> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=7985 $D=0
M85 WL<48> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=9520 $D=0
M86 WL<47> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=11475 $D=0
M87 WL<46> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=13010 $D=0
M88 WL<45> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=14545 $D=0
M89 WL<44> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=16080 $D=0
M90 WL<43> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=17615 $D=0
M91 WL<42> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=19150 $D=0
M92 WL<41> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=20685 $D=0
M93 WL<40> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=22220 $D=0
M94 WL<39> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=23755 $D=0
M95 WL<38> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=25290 $D=0
M96 WL<37> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=26825 $D=0
M97 WL<36> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=28360 $D=0
M98 WL<35> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=29895 $D=0
M99 WL<34> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=31430 $D=0
M100 WL<33> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=32965 $D=0
M101 WL<32> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=34500 $D=0
M102 WL<31> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=36455 $D=0
M103 WL<30> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=37990 $D=0
M104 WL<29> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=39525 $D=0
M105 WL<28> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=41060 $D=0
M106 WL<27> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=42595 $D=0
M107 WL<26> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=44130 $D=0
M108 WL<25> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=45665 $D=0
M109 WL<24> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=47200 $D=0
M110 WL<23> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=48735 $D=0
M111 WL<22> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=50270 $D=0
M112 WL<21> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=51805 $D=0
M113 WL<20> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=53340 $D=0
M114 WL<19> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=54875 $D=0
M115 WL<18> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=56410 $D=0
M116 WL<17> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=57945 $D=0
M117 WL<16> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=59480 $D=0
M118 WL<15> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=61435 $D=0
M119 WL<14> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=62970 $D=0
M120 WL<13> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=64505 $D=0
M121 WL<12> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=66040 $D=0
M122 WL<11> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=67575 $D=0
M123 WL<10> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=69110 $D=0
M124 WL<9> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=70645 $D=0
M125 WL<8> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=72180 $D=0
M126 WL<7> 24 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=73715 $D=0
M127 WL<6> 25 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=75250 $D=0
M128 WL<5> 26 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=76785 $D=0
M129 WL<4> 27 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=78320 $D=0
M130 WL<3> 28 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=79855 $D=0
M131 WL<2> 29 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=81390 $D=0
M132 WL<1> 30 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=82925 $D=0
M133 WL<0> 31 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-40590 $Y=84460 $D=0
M134 WL<63> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-13505 $D=0
M135 WL<62> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-11970 $D=0
M136 WL<61> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-10435 $D=0
M137 WL<60> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-8900 $D=0
M138 WL<59> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-7365 $D=0
M139 WL<58> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-5830 $D=0
M140 WL<57> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-4295 $D=0
M141 WL<56> 16 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-2760 $D=0
M142 WL<55> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=-1225 $D=0
M143 WL<54> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=310 $D=0
M144 WL<53> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=1845 $D=0
M145 WL<52> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=3380 $D=0
M146 WL<51> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=4915 $D=0
M147 WL<50> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=6450 $D=0
M148 WL<49> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=7985 $D=0
M149 WL<48> 17 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=9520 $D=0
M150 WL<47> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=11475 $D=0
M151 WL<46> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=13010 $D=0
M152 WL<45> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=14545 $D=0
M153 WL<44> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=16080 $D=0
M154 WL<43> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=17615 $D=0
M155 WL<42> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=19150 $D=0
M156 WL<41> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=20685 $D=0
M157 WL<40> 18 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=22220 $D=0
M158 WL<39> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=23755 $D=0
M159 WL<38> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=25290 $D=0
M160 WL<37> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=26825 $D=0
M161 WL<36> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=28360 $D=0
M162 WL<35> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=29895 $D=0
M163 WL<34> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=31430 $D=0
M164 WL<33> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=32965 $D=0
M165 WL<32> 19 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=34500 $D=0
M166 WL<31> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=36455 $D=0
M167 WL<30> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=37990 $D=0
M168 WL<29> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=39525 $D=0
M169 WL<28> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=41060 $D=0
M170 WL<27> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=42595 $D=0
M171 WL<26> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=44130 $D=0
M172 WL<25> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=45665 $D=0
M173 WL<24> 20 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=47200 $D=0
M174 WL<23> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=48735 $D=0
M175 WL<22> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=50270 $D=0
M176 WL<21> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=51805 $D=0
M177 WL<20> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=53340 $D=0
M178 WL<19> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=54875 $D=0
M179 WL<18> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=56410 $D=0
M180 WL<17> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=57945 $D=0
M181 WL<16> 21 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=59480 $D=0
M182 WL<15> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=61435 $D=0
M183 WL<14> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=62970 $D=0
M184 WL<13> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=64505 $D=0
M185 WL<12> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=66040 $D=0
M186 WL<11> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=67575 $D=0
M187 WL<10> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=69110 $D=0
M188 WL<9> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=70645 $D=0
M189 WL<8> 22 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=72180 $D=0
M190 WL<7> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=73715 $D=0
M191 WL<6> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=75250 $D=0
M192 WL<5> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=76785 $D=0
M193 WL<4> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=78320 $D=0
M194 WL<3> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=79855 $D=0
M195 WL<2> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=81390 $D=0
M196 WL<1> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=82925 $D=0
M197 WL<0> 23 VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-39440 $Y=84460 $D=0
M198 VSS WL<63> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-13645 $D=0
M199 VSS WL<62> 263 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-12110 $D=0
M200 VSS WL<61> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-10575 $D=0
M201 VSS WL<60> 264 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-9040 $D=0
M202 VSS WL<59> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-7505 $D=0
M203 VSS WL<58> 265 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-5970 $D=0
M204 VSS WL<57> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-4435 $D=0
M205 VSS WL<56> 266 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-2900 $D=0
M206 VSS WL<55> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=-1365 $D=0
M207 VSS WL<54> 267 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=170 $D=0
M208 VSS WL<53> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=1705 $D=0
M209 VSS WL<52> 268 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=3240 $D=0
M210 VSS WL<51> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=4775 $D=0
M211 VSS WL<50> 269 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=6310 $D=0
M212 VSS WL<49> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=7845 $D=0
M213 VSS WL<48> 270 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=9380 $D=0
M214 VSS WL<47> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=11335 $D=0
M215 VSS WL<46> 271 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=12870 $D=0
M216 VSS WL<45> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=14405 $D=0
M217 VSS WL<44> 272 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=15940 $D=0
M218 VSS WL<43> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=17475 $D=0
M219 VSS WL<42> 273 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=19010 $D=0
M220 VSS WL<41> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=20545 $D=0
M221 VSS WL<40> 274 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=22080 $D=0
M222 VSS WL<39> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=23615 $D=0
M223 VSS WL<38> 275 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=25150 $D=0
M224 VSS WL<37> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=26685 $D=0
M225 VSS WL<36> 276 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=28220 $D=0
M226 VSS WL<35> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=29755 $D=0
M227 VSS WL<34> 277 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=31290 $D=0
M228 VSS WL<33> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=32825 $D=0
M229 VSS WL<32> 278 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=34360 $D=0
M230 VSS WL<31> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=36315 $D=0
M231 VSS WL<30> 279 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=37850 $D=0
M232 VSS WL<29> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=39385 $D=0
M233 VSS WL<28> 280 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=40920 $D=0
M234 VSS WL<27> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=42455 $D=0
M235 VSS WL<26> 281 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=43990 $D=0
M236 VSS WL<25> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=45525 $D=0
M237 VSS WL<24> 282 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=47060 $D=0
M238 VSS WL<23> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=48595 $D=0
M239 VSS WL<22> 283 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=50130 $D=0
M240 VSS WL<21> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=51665 $D=0
M241 VSS WL<20> 284 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=53200 $D=0
M242 VSS WL<19> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=54735 $D=0
M243 VSS WL<18> 285 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=56270 $D=0
M244 VSS WL<17> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=57805 $D=0
M245 VSS WL<16> 286 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=59340 $D=0
M246 VSS WL<15> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=61295 $D=0
M247 VSS WL<14> 287 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=62830 $D=0
M248 VSS WL<13> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=64365 $D=0
M249 VSS WL<12> 288 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=65900 $D=0
M250 VSS WL<11> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=67435 $D=0
M251 VSS WL<10> 289 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=68970 $D=0
M252 VSS WL<9> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=70505 $D=0
M253 VSS WL<8> 290 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=72040 $D=0
M254 VSS WL<7> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=73575 $D=0
M255 VSS WL<6> 291 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=75110 $D=0
M256 VSS WL<5> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=76645 $D=0
M257 VSS WL<4> 292 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=78180 $D=0
M258 VSS WL<3> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=79715 $D=0
M259 VSS WL<2> 293 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=81250 $D=0
M260 VSS WL<1> BL<0> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=82785 $D=0
M261 VSS WL<0> 294 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-27660 $Y=84320 $D=0
M262 130 YOUT<1> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27314 $Y=-35070 $D=0
M263 131 YOUT<0> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27314 $Y=-25360 $D=0
M264 BL<1> YOUT<1> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27129 $Y=-37036 $D=0
M265 BL<0> YOUT<0> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-27129 $Y=-27326 $D=0
M266 295 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-13645 $D=0
M267 BL<1> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-12110 $D=0
M268 296 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-10575 $D=0
M269 BL<1> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-9040 $D=0
M270 297 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-7505 $D=0
M271 BL<1> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-5970 $D=0
M272 298 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-4435 $D=0
M273 BL<1> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-2900 $D=0
M274 299 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=-1365 $D=0
M275 BL<1> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=170 $D=0
M276 300 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=1705 $D=0
M277 BL<1> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=3240 $D=0
M278 301 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=4775 $D=0
M279 BL<1> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=6310 $D=0
M280 302 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=7845 $D=0
M281 BL<1> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=9380 $D=0
M282 303 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=11335 $D=0
M283 BL<1> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=12870 $D=0
M284 304 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=14405 $D=0
M285 BL<1> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=15940 $D=0
M286 305 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=17475 $D=0
M287 BL<1> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=19010 $D=0
M288 306 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=20545 $D=0
M289 BL<1> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=22080 $D=0
M290 307 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=23615 $D=0
M291 BL<1> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=25150 $D=0
M292 308 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=26685 $D=0
M293 BL<1> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=28220 $D=0
M294 309 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=29755 $D=0
M295 BL<1> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=31290 $D=0
M296 310 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=32825 $D=0
M297 BL<1> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=34360 $D=0
M298 311 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=36315 $D=0
M299 BL<1> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=37850 $D=0
M300 312 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=39385 $D=0
M301 BL<1> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=40920 $D=0
M302 313 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=42455 $D=0
M303 BL<1> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=43990 $D=0
M304 314 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=45525 $D=0
M305 BL<1> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=47060 $D=0
M306 315 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=48595 $D=0
M307 BL<1> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=50130 $D=0
M308 316 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=51665 $D=0
M309 BL<1> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=53200 $D=0
M310 317 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=54735 $D=0
M311 BL<1> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=56270 $D=0
M312 318 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=57805 $D=0
M313 BL<1> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=59340 $D=0
M314 319 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=61295 $D=0
M315 BL<1> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=62830 $D=0
M316 320 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=64365 $D=0
M317 BL<1> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=65900 $D=0
M318 321 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=67435 $D=0
M319 BL<1> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=68970 $D=0
M320 322 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=70505 $D=0
M321 BL<1> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=72040 $D=0
M322 323 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=73575 $D=0
M323 BL<1> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=75110 $D=0
M324 324 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=76645 $D=0
M325 BL<1> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=78180 $D=0
M326 325 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=79715 $D=0
M327 BL<1> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=81250 $D=0
M328 326 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=82785 $D=0
M329 BL<1> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-26970 $Y=84320 $D=0
M330 VSS WL<63> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-13645 $D=0
M331 VSS WL<62> 327 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-12110 $D=0
M332 VSS WL<61> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-10575 $D=0
M333 VSS WL<60> 328 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-9040 $D=0
M334 VSS WL<59> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-7505 $D=0
M335 VSS WL<58> 329 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-5970 $D=0
M336 VSS WL<57> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-4435 $D=0
M337 VSS WL<56> 330 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-2900 $D=0
M338 VSS WL<55> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=-1365 $D=0
M339 VSS WL<54> 331 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=170 $D=0
M340 VSS WL<53> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=1705 $D=0
M341 VSS WL<52> 332 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=3240 $D=0
M342 VSS WL<51> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=4775 $D=0
M343 VSS WL<50> 333 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=6310 $D=0
M344 VSS WL<49> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=7845 $D=0
M345 VSS WL<48> 334 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=9380 $D=0
M346 VSS WL<47> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=11335 $D=0
M347 VSS WL<46> 335 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=12870 $D=0
M348 VSS WL<45> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=14405 $D=0
M349 VSS WL<44> 336 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=15940 $D=0
M350 VSS WL<43> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=17475 $D=0
M351 VSS WL<42> 337 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=19010 $D=0
M352 VSS WL<41> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=20545 $D=0
M353 VSS WL<40> 338 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=22080 $D=0
M354 VSS WL<39> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=23615 $D=0
M355 VSS WL<38> 339 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=25150 $D=0
M356 VSS WL<37> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=26685 $D=0
M357 VSS WL<36> 340 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=28220 $D=0
M358 VSS WL<35> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=29755 $D=0
M359 VSS WL<34> 341 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=31290 $D=0
M360 VSS WL<33> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=32825 $D=0
M361 VSS WL<32> 342 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=34360 $D=0
M362 VSS WL<31> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=36315 $D=0
M363 VSS WL<30> 343 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=37850 $D=0
M364 VSS WL<29> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=39385 $D=0
M365 VSS WL<28> 344 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=40920 $D=0
M366 VSS WL<27> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=42455 $D=0
M367 VSS WL<26> 345 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=43990 $D=0
M368 VSS WL<25> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=45525 $D=0
M369 VSS WL<24> 346 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=47060 $D=0
M370 VSS WL<23> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=48595 $D=0
M371 VSS WL<22> 347 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=50130 $D=0
M372 VSS WL<21> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=51665 $D=0
M373 VSS WL<20> 348 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=53200 $D=0
M374 VSS WL<19> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=54735 $D=0
M375 VSS WL<18> 349 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=56270 $D=0
M376 VSS WL<17> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=57805 $D=0
M377 VSS WL<16> 350 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=59340 $D=0
M378 VSS WL<15> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=61295 $D=0
M379 VSS WL<14> 351 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=62830 $D=0
M380 VSS WL<13> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=64365 $D=0
M381 VSS WL<12> 352 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=65900 $D=0
M382 VSS WL<11> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=67435 $D=0
M383 VSS WL<10> 353 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=68970 $D=0
M384 VSS WL<9> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=70505 $D=0
M385 VSS WL<8> 354 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=72040 $D=0
M386 VSS WL<7> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=73575 $D=0
M387 VSS WL<6> 355 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=75110 $D=0
M388 VSS WL<5> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=76645 $D=0
M389 VSS WL<4> 356 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=78180 $D=0
M390 VSS WL<3> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=79715 $D=0
M391 VSS WL<2> 357 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=81250 $D=0
M392 VSS WL<1> BL<2> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=82785 $D=0
M393 VSS WL<0> 358 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-25510 $Y=84320 $D=0
M394 132 YOUT<3> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-25164 $Y=-35070 $D=0
M395 133 YOUT<2> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-25164 $Y=-25360 $D=0
M396 BL<3> YOUT<3> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-24979 $Y=-37036 $D=0
M397 BL<2> YOUT<2> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-24979 $Y=-27326 $D=0
M398 359 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-13645 $D=0
M399 BL<3> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-12110 $D=0
M400 360 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-10575 $D=0
M401 BL<3> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-9040 $D=0
M402 361 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-7505 $D=0
M403 BL<3> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-5970 $D=0
M404 362 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-4435 $D=0
M405 BL<3> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-2900 $D=0
M406 363 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=-1365 $D=0
M407 BL<3> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=170 $D=0
M408 364 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=1705 $D=0
M409 BL<3> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=3240 $D=0
M410 365 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=4775 $D=0
M411 BL<3> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=6310 $D=0
M412 366 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=7845 $D=0
M413 BL<3> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=9380 $D=0
M414 367 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=11335 $D=0
M415 BL<3> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=12870 $D=0
M416 368 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=14405 $D=0
M417 BL<3> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=15940 $D=0
M418 369 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=17475 $D=0
M419 BL<3> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=19010 $D=0
M420 370 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=20545 $D=0
M421 BL<3> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=22080 $D=0
M422 371 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=23615 $D=0
M423 BL<3> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=25150 $D=0
M424 372 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=26685 $D=0
M425 BL<3> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=28220 $D=0
M426 373 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=29755 $D=0
M427 BL<3> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=31290 $D=0
M428 374 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=32825 $D=0
M429 BL<3> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=34360 $D=0
M430 375 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=36315 $D=0
M431 BL<3> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=37850 $D=0
M432 376 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=39385 $D=0
M433 BL<3> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=40920 $D=0
M434 377 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=42455 $D=0
M435 BL<3> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=43990 $D=0
M436 378 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=45525 $D=0
M437 BL<3> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=47060 $D=0
M438 379 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=48595 $D=0
M439 BL<3> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=50130 $D=0
M440 380 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=51665 $D=0
M441 BL<3> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=53200 $D=0
M442 381 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=54735 $D=0
M443 BL<3> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=56270 $D=0
M444 382 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=57805 $D=0
M445 BL<3> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=59340 $D=0
M446 383 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=61295 $D=0
M447 BL<3> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=62830 $D=0
M448 384 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=64365 $D=0
M449 BL<3> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=65900 $D=0
M450 385 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=67435 $D=0
M451 BL<3> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=68970 $D=0
M452 386 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=70505 $D=0
M453 BL<3> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=72040 $D=0
M454 387 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=73575 $D=0
M455 BL<3> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=75110 $D=0
M456 388 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=76645 $D=0
M457 BL<3> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=78180 $D=0
M458 389 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=79715 $D=0
M459 BL<3> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=81250 $D=0
M460 390 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=82785 $D=0
M461 BL<3> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-24820 $Y=84320 $D=0
M462 VSS WL<63> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-13645 $D=0
M463 VSS WL<62> 391 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-12110 $D=0
M464 VSS WL<61> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-10575 $D=0
M465 VSS WL<60> 392 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-9040 $D=0
M466 VSS WL<59> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-7505 $D=0
M467 VSS WL<58> 393 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-5970 $D=0
M468 VSS WL<57> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-4435 $D=0
M469 VSS WL<56> 394 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-2900 $D=0
M470 VSS WL<55> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=-1365 $D=0
M471 VSS WL<54> 395 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=170 $D=0
M472 VSS WL<53> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=1705 $D=0
M473 VSS WL<52> 396 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=3240 $D=0
M474 VSS WL<51> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=4775 $D=0
M475 VSS WL<50> 397 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=6310 $D=0
M476 VSS WL<49> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=7845 $D=0
M477 VSS WL<48> 398 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=9380 $D=0
M478 VSS WL<47> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=11335 $D=0
M479 VSS WL<46> 399 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=12870 $D=0
M480 VSS WL<45> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=14405 $D=0
M481 VSS WL<44> 400 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=15940 $D=0
M482 VSS WL<43> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=17475 $D=0
M483 VSS WL<42> 401 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=19010 $D=0
M484 VSS WL<41> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=20545 $D=0
M485 VSS WL<40> 402 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=22080 $D=0
M486 VSS WL<39> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=23615 $D=0
M487 VSS WL<38> 403 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=25150 $D=0
M488 VSS WL<37> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=26685 $D=0
M489 VSS WL<36> 404 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=28220 $D=0
M490 VSS WL<35> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=29755 $D=0
M491 VSS WL<34> 405 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=31290 $D=0
M492 VSS WL<33> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=32825 $D=0
M493 VSS WL<32> 406 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=34360 $D=0
M494 VSS WL<31> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=36315 $D=0
M495 VSS WL<30> 407 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=37850 $D=0
M496 VSS WL<29> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=39385 $D=0
M497 VSS WL<28> 408 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=40920 $D=0
M498 VSS WL<27> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=42455 $D=0
M499 VSS WL<26> 409 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=43990 $D=0
M500 VSS WL<25> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=45525 $D=0
M501 VSS WL<24> 410 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=47060 $D=0
M502 VSS WL<23> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=48595 $D=0
M503 VSS WL<22> 411 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=50130 $D=0
M504 VSS WL<21> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=51665 $D=0
M505 VSS WL<20> 412 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=53200 $D=0
M506 VSS WL<19> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=54735 $D=0
M507 VSS WL<18> 413 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=56270 $D=0
M508 VSS WL<17> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=57805 $D=0
M509 VSS WL<16> 414 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=59340 $D=0
M510 VSS WL<15> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=61295 $D=0
M511 VSS WL<14> 415 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=62830 $D=0
M512 VSS WL<13> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=64365 $D=0
M513 VSS WL<12> 416 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=65900 $D=0
M514 VSS WL<11> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=67435 $D=0
M515 VSS WL<10> 417 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=68970 $D=0
M516 VSS WL<9> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=70505 $D=0
M517 VSS WL<8> 418 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=72040 $D=0
M518 VSS WL<7> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=73575 $D=0
M519 VSS WL<6> 419 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=75110 $D=0
M520 VSS WL<5> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=76645 $D=0
M521 VSS WL<4> 420 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=78180 $D=0
M522 VSS WL<3> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=79715 $D=0
M523 VSS WL<2> 421 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=81250 $D=0
M524 VSS WL<1> BL<4> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=82785 $D=0
M525 VSS WL<0> 422 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-23360 $Y=84320 $D=0
M526 134 YOUT<5> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-23014 $Y=-35070 $D=0
M527 135 YOUT<4> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-23014 $Y=-25360 $D=0
M528 BL<5> YOUT<5> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-22829 $Y=-37036 $D=0
M529 BL<4> YOUT<4> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-22829 $Y=-27326 $D=0
M530 423 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-13645 $D=0
M531 BL<5> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-12110 $D=0
M532 424 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-10575 $D=0
M533 BL<5> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-9040 $D=0
M534 425 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-7505 $D=0
M535 BL<5> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-5970 $D=0
M536 426 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-4435 $D=0
M537 BL<5> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-2900 $D=0
M538 427 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=-1365 $D=0
M539 BL<5> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=170 $D=0
M540 428 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=1705 $D=0
M541 BL<5> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=3240 $D=0
M542 429 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=4775 $D=0
M543 BL<5> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=6310 $D=0
M544 430 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=7845 $D=0
M545 BL<5> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=9380 $D=0
M546 431 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=11335 $D=0
M547 BL<5> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=12870 $D=0
M548 432 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=14405 $D=0
M549 BL<5> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=15940 $D=0
M550 433 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=17475 $D=0
M551 BL<5> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=19010 $D=0
M552 434 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=20545 $D=0
M553 BL<5> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=22080 $D=0
M554 435 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=23615 $D=0
M555 BL<5> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=25150 $D=0
M556 436 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=26685 $D=0
M557 BL<5> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=28220 $D=0
M558 437 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=29755 $D=0
M559 BL<5> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=31290 $D=0
M560 438 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=32825 $D=0
M561 BL<5> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=34360 $D=0
M562 439 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=36315 $D=0
M563 BL<5> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=37850 $D=0
M564 440 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=39385 $D=0
M565 BL<5> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=40920 $D=0
M566 441 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=42455 $D=0
M567 BL<5> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=43990 $D=0
M568 442 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=45525 $D=0
M569 BL<5> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=47060 $D=0
M570 443 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=48595 $D=0
M571 BL<5> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=50130 $D=0
M572 444 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=51665 $D=0
M573 BL<5> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=53200 $D=0
M574 445 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=54735 $D=0
M575 BL<5> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=56270 $D=0
M576 446 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=57805 $D=0
M577 BL<5> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=59340 $D=0
M578 447 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=61295 $D=0
M579 BL<5> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=62830 $D=0
M580 448 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=64365 $D=0
M581 BL<5> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=65900 $D=0
M582 449 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=67435 $D=0
M583 BL<5> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=68970 $D=0
M584 450 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=70505 $D=0
M585 BL<5> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=72040 $D=0
M586 451 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=73575 $D=0
M587 BL<5> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=75110 $D=0
M588 452 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=76645 $D=0
M589 BL<5> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=78180 $D=0
M590 453 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=79715 $D=0
M591 BL<5> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=81250 $D=0
M592 454 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=82785 $D=0
M593 BL<5> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-22670 $Y=84320 $D=0
M594 VSS WL<63> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-13645 $D=0
M595 VSS WL<62> 455 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-12110 $D=0
M596 VSS WL<61> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-10575 $D=0
M597 VSS WL<60> 456 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-9040 $D=0
M598 VSS WL<59> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-7505 $D=0
M599 VSS WL<58> 457 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-5970 $D=0
M600 VSS WL<57> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-4435 $D=0
M601 VSS WL<56> 458 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-2900 $D=0
M602 VSS WL<55> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=-1365 $D=0
M603 VSS WL<54> 459 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=170 $D=0
M604 VSS WL<53> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=1705 $D=0
M605 VSS WL<52> 460 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=3240 $D=0
M606 VSS WL<51> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=4775 $D=0
M607 VSS WL<50> 461 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=6310 $D=0
M608 VSS WL<49> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=7845 $D=0
M609 VSS WL<48> 462 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=9380 $D=0
M610 VSS WL<47> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=11335 $D=0
M611 VSS WL<46> 463 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=12870 $D=0
M612 VSS WL<45> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=14405 $D=0
M613 VSS WL<44> 464 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=15940 $D=0
M614 VSS WL<43> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=17475 $D=0
M615 VSS WL<42> 465 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=19010 $D=0
M616 VSS WL<41> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=20545 $D=0
M617 VSS WL<40> 466 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=22080 $D=0
M618 VSS WL<39> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=23615 $D=0
M619 VSS WL<38> 467 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=25150 $D=0
M620 VSS WL<37> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=26685 $D=0
M621 VSS WL<36> 468 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=28220 $D=0
M622 VSS WL<35> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=29755 $D=0
M623 VSS WL<34> 469 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=31290 $D=0
M624 VSS WL<33> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=32825 $D=0
M625 VSS WL<32> 470 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=34360 $D=0
M626 VSS WL<31> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=36315 $D=0
M627 VSS WL<30> 471 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=37850 $D=0
M628 VSS WL<29> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=39385 $D=0
M629 VSS WL<28> 472 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=40920 $D=0
M630 VSS WL<27> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=42455 $D=0
M631 VSS WL<26> 473 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=43990 $D=0
M632 VSS WL<25> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=45525 $D=0
M633 VSS WL<24> 474 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=47060 $D=0
M634 VSS WL<23> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=48595 $D=0
M635 VSS WL<22> 475 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=50130 $D=0
M636 VSS WL<21> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=51665 $D=0
M637 VSS WL<20> 476 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=53200 $D=0
M638 VSS WL<19> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=54735 $D=0
M639 VSS WL<18> 477 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=56270 $D=0
M640 VSS WL<17> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=57805 $D=0
M641 VSS WL<16> 478 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=59340 $D=0
M642 VSS WL<15> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=61295 $D=0
M643 VSS WL<14> 479 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=62830 $D=0
M644 VSS WL<13> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=64365 $D=0
M645 VSS WL<12> 480 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=65900 $D=0
M646 VSS WL<11> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=67435 $D=0
M647 VSS WL<10> 481 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=68970 $D=0
M648 VSS WL<9> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=70505 $D=0
M649 VSS WL<8> 482 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=72040 $D=0
M650 VSS WL<7> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=73575 $D=0
M651 VSS WL<6> 483 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=75110 $D=0
M652 VSS WL<5> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=76645 $D=0
M653 VSS WL<4> 484 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=78180 $D=0
M654 VSS WL<3> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=79715 $D=0
M655 VSS WL<2> 485 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=81250 $D=0
M656 VSS WL<1> BL<6> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=82785 $D=0
M657 VSS WL<0> 486 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-21210 $Y=84320 $D=0
M658 136 YOUT<7> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20864 $Y=-35070 $D=0
M659 137 YOUT<6> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20864 $Y=-25360 $D=0
M660 BL<7> YOUT<7> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20679 $Y=-37036 $D=0
M661 BL<6> YOUT<6> DL<0> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-20679 $Y=-27326 $D=0
M662 487 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-13645 $D=0
M663 BL<7> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-12110 $D=0
M664 488 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-10575 $D=0
M665 BL<7> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-9040 $D=0
M666 489 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-7505 $D=0
M667 BL<7> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-5970 $D=0
M668 490 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-4435 $D=0
M669 BL<7> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-2900 $D=0
M670 491 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=-1365 $D=0
M671 BL<7> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=170 $D=0
M672 492 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=1705 $D=0
M673 BL<7> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=3240 $D=0
M674 493 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=4775 $D=0
M675 BL<7> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=6310 $D=0
M676 494 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=7845 $D=0
M677 BL<7> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=9380 $D=0
M678 495 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=11335 $D=0
M679 BL<7> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=12870 $D=0
M680 496 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=14405 $D=0
M681 BL<7> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=15940 $D=0
M682 497 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=17475 $D=0
M683 BL<7> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=19010 $D=0
M684 498 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=20545 $D=0
M685 BL<7> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=22080 $D=0
M686 499 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=23615 $D=0
M687 BL<7> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=25150 $D=0
M688 500 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=26685 $D=0
M689 BL<7> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=28220 $D=0
M690 501 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=29755 $D=0
M691 BL<7> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=31290 $D=0
M692 502 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=32825 $D=0
M693 BL<7> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=34360 $D=0
M694 503 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=36315 $D=0
M695 BL<7> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=37850 $D=0
M696 504 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=39385 $D=0
M697 BL<7> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=40920 $D=0
M698 505 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=42455 $D=0
M699 BL<7> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=43990 $D=0
M700 506 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=45525 $D=0
M701 BL<7> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=47060 $D=0
M702 507 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=48595 $D=0
M703 BL<7> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=50130 $D=0
M704 508 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=51665 $D=0
M705 BL<7> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=53200 $D=0
M706 509 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=54735 $D=0
M707 BL<7> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=56270 $D=0
M708 510 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=57805 $D=0
M709 BL<7> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=59340 $D=0
M710 511 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=61295 $D=0
M711 BL<7> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=62830 $D=0
M712 512 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=64365 $D=0
M713 BL<7> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=65900 $D=0
M714 513 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=67435 $D=0
M715 BL<7> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=68970 $D=0
M716 514 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=70505 $D=0
M717 BL<7> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=72040 $D=0
M718 515 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=73575 $D=0
M719 BL<7> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=75110 $D=0
M720 516 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=76645 $D=0
M721 BL<7> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=78180 $D=0
M722 517 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=79715 $D=0
M723 BL<7> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=81250 $D=0
M724 518 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=82785 $D=0
M725 BL<7> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-20520 $Y=84320 $D=0
M726 VSS WL<63> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-13645 $D=0
M727 VSS WL<62> 519 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-12110 $D=0
M728 VSS WL<61> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-10575 $D=0
M729 VSS WL<60> 520 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-9040 $D=0
M730 VSS WL<59> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-7505 $D=0
M731 VSS WL<58> 521 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-5970 $D=0
M732 VSS WL<57> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-4435 $D=0
M733 VSS WL<56> 522 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-2900 $D=0
M734 VSS WL<55> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=-1365 $D=0
M735 VSS WL<54> 523 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=170 $D=0
M736 VSS WL<53> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=1705 $D=0
M737 VSS WL<52> 524 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=3240 $D=0
M738 VSS WL<51> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=4775 $D=0
M739 VSS WL<50> 525 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=6310 $D=0
M740 VSS WL<49> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=7845 $D=0
M741 VSS WL<48> 526 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=9380 $D=0
M742 VSS WL<47> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=11335 $D=0
M743 VSS WL<46> 527 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=12870 $D=0
M744 VSS WL<45> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=14405 $D=0
M745 VSS WL<44> 528 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=15940 $D=0
M746 VSS WL<43> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=17475 $D=0
M747 VSS WL<42> 529 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=19010 $D=0
M748 VSS WL<41> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=20545 $D=0
M749 VSS WL<40> 530 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=22080 $D=0
M750 VSS WL<39> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=23615 $D=0
M751 VSS WL<38> 531 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=25150 $D=0
M752 VSS WL<37> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=26685 $D=0
M753 VSS WL<36> 532 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=28220 $D=0
M754 VSS WL<35> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=29755 $D=0
M755 VSS WL<34> 533 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=31290 $D=0
M756 VSS WL<33> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=32825 $D=0
M757 VSS WL<32> 534 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=34360 $D=0
M758 VSS WL<31> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=36315 $D=0
M759 VSS WL<30> 535 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=37850 $D=0
M760 VSS WL<29> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=39385 $D=0
M761 VSS WL<28> 536 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=40920 $D=0
M762 VSS WL<27> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=42455 $D=0
M763 VSS WL<26> 537 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=43990 $D=0
M764 VSS WL<25> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=45525 $D=0
M765 VSS WL<24> 538 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=47060 $D=0
M766 VSS WL<23> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=48595 $D=0
M767 VSS WL<22> 539 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=50130 $D=0
M768 VSS WL<21> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=51665 $D=0
M769 VSS WL<20> 540 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=53200 $D=0
M770 VSS WL<19> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=54735 $D=0
M771 VSS WL<18> 541 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=56270 $D=0
M772 VSS WL<17> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=57805 $D=0
M773 VSS WL<16> 542 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=59340 $D=0
M774 VSS WL<15> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=61295 $D=0
M775 VSS WL<14> 543 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=62830 $D=0
M776 VSS WL<13> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=64365 $D=0
M777 VSS WL<12> 544 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=65900 $D=0
M778 VSS WL<11> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=67435 $D=0
M779 VSS WL<10> 545 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=68970 $D=0
M780 VSS WL<9> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=70505 $D=0
M781 VSS WL<8> 546 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=72040 $D=0
M782 VSS WL<7> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=73575 $D=0
M783 VSS WL<6> 547 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=75110 $D=0
M784 VSS WL<5> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=76645 $D=0
M785 VSS WL<4> 548 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=78180 $D=0
M786 VSS WL<3> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=79715 $D=0
M787 VSS WL<2> 549 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=81250 $D=0
M788 VSS WL<1> BL<8> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=82785 $D=0
M789 VSS WL<0> 550 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-19060 $Y=84320 $D=0
M790 138 YOUT<1> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18714 $Y=-35070 $D=0
M791 139 YOUT<0> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18714 $Y=-25360 $D=0
M792 BL<9> YOUT<1> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18529 $Y=-37036 $D=0
M793 BL<8> YOUT<0> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-18529 $Y=-27326 $D=0
M794 551 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-13645 $D=0
M795 BL<9> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-12110 $D=0
M796 552 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-10575 $D=0
M797 BL<9> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-9040 $D=0
M798 553 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-7505 $D=0
M799 BL<9> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-5970 $D=0
M800 554 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-4435 $D=0
M801 BL<9> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-2900 $D=0
M802 555 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=-1365 $D=0
M803 BL<9> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=170 $D=0
M804 556 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=1705 $D=0
M805 BL<9> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=3240 $D=0
M806 557 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=4775 $D=0
M807 BL<9> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=6310 $D=0
M808 558 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=7845 $D=0
M809 BL<9> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=9380 $D=0
M810 559 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=11335 $D=0
M811 BL<9> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=12870 $D=0
M812 560 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=14405 $D=0
M813 BL<9> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=15940 $D=0
M814 561 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=17475 $D=0
M815 BL<9> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=19010 $D=0
M816 562 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=20545 $D=0
M817 BL<9> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=22080 $D=0
M818 563 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=23615 $D=0
M819 BL<9> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=25150 $D=0
M820 564 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=26685 $D=0
M821 BL<9> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=28220 $D=0
M822 565 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=29755 $D=0
M823 BL<9> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=31290 $D=0
M824 566 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=32825 $D=0
M825 BL<9> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=34360 $D=0
M826 567 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=36315 $D=0
M827 BL<9> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=37850 $D=0
M828 568 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=39385 $D=0
M829 BL<9> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=40920 $D=0
M830 569 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=42455 $D=0
M831 BL<9> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=43990 $D=0
M832 570 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=45525 $D=0
M833 BL<9> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=47060 $D=0
M834 571 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=48595 $D=0
M835 BL<9> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=50130 $D=0
M836 572 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=51665 $D=0
M837 BL<9> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=53200 $D=0
M838 573 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=54735 $D=0
M839 BL<9> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=56270 $D=0
M840 574 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=57805 $D=0
M841 BL<9> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=59340 $D=0
M842 575 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=61295 $D=0
M843 BL<9> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=62830 $D=0
M844 576 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=64365 $D=0
M845 BL<9> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=65900 $D=0
M846 577 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=67435 $D=0
M847 BL<9> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=68970 $D=0
M848 578 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=70505 $D=0
M849 BL<9> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=72040 $D=0
M850 579 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=73575 $D=0
M851 BL<9> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=75110 $D=0
M852 580 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=76645 $D=0
M853 BL<9> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=78180 $D=0
M854 581 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=79715 $D=0
M855 BL<9> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=81250 $D=0
M856 582 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=82785 $D=0
M857 BL<9> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-18370 $Y=84320 $D=0
M858 VSS WL<63> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-13645 $D=0
M859 VSS WL<62> 583 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-12110 $D=0
M860 VSS WL<61> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-10575 $D=0
M861 VSS WL<60> 584 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-9040 $D=0
M862 VSS WL<59> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-7505 $D=0
M863 VSS WL<58> 585 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-5970 $D=0
M864 VSS WL<57> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-4435 $D=0
M865 VSS WL<56> 586 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-2900 $D=0
M866 VSS WL<55> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=-1365 $D=0
M867 VSS WL<54> 587 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=170 $D=0
M868 VSS WL<53> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=1705 $D=0
M869 VSS WL<52> 588 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=3240 $D=0
M870 VSS WL<51> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=4775 $D=0
M871 VSS WL<50> 589 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=6310 $D=0
M872 VSS WL<49> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=7845 $D=0
M873 VSS WL<48> 590 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=9380 $D=0
M874 VSS WL<47> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=11335 $D=0
M875 VSS WL<46> 591 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=12870 $D=0
M876 VSS WL<45> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=14405 $D=0
M877 VSS WL<44> 592 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=15940 $D=0
M878 VSS WL<43> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=17475 $D=0
M879 VSS WL<42> 593 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=19010 $D=0
M880 VSS WL<41> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=20545 $D=0
M881 VSS WL<40> 594 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=22080 $D=0
M882 VSS WL<39> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=23615 $D=0
M883 VSS WL<38> 595 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=25150 $D=0
M884 VSS WL<37> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=26685 $D=0
M885 VSS WL<36> 596 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=28220 $D=0
M886 VSS WL<35> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=29755 $D=0
M887 VSS WL<34> 597 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=31290 $D=0
M888 VSS WL<33> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=32825 $D=0
M889 VSS WL<32> 598 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=34360 $D=0
M890 VSS WL<31> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=36315 $D=0
M891 VSS WL<30> 599 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=37850 $D=0
M892 VSS WL<29> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=39385 $D=0
M893 VSS WL<28> 600 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=40920 $D=0
M894 VSS WL<27> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=42455 $D=0
M895 VSS WL<26> 601 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=43990 $D=0
M896 VSS WL<25> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=45525 $D=0
M897 VSS WL<24> 602 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=47060 $D=0
M898 VSS WL<23> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=48595 $D=0
M899 VSS WL<22> 603 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=50130 $D=0
M900 VSS WL<21> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=51665 $D=0
M901 VSS WL<20> 604 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=53200 $D=0
M902 VSS WL<19> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=54735 $D=0
M903 VSS WL<18> 605 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=56270 $D=0
M904 VSS WL<17> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=57805 $D=0
M905 VSS WL<16> 606 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=59340 $D=0
M906 VSS WL<15> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=61295 $D=0
M907 VSS WL<14> 607 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=62830 $D=0
M908 VSS WL<13> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=64365 $D=0
M909 VSS WL<12> 608 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=65900 $D=0
M910 VSS WL<11> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=67435 $D=0
M911 VSS WL<10> 609 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=68970 $D=0
M912 VSS WL<9> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=70505 $D=0
M913 VSS WL<8> 610 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=72040 $D=0
M914 VSS WL<7> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=73575 $D=0
M915 VSS WL<6> 611 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=75110 $D=0
M916 VSS WL<5> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=76645 $D=0
M917 VSS WL<4> 612 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=78180 $D=0
M918 VSS WL<3> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=79715 $D=0
M919 VSS WL<2> 613 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=81250 $D=0
M920 VSS WL<1> BL<10> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=82785 $D=0
M921 VSS WL<0> 614 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-16910 $Y=84320 $D=0
M922 140 YOUT<3> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16564 $Y=-35070 $D=0
M923 141 YOUT<2> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16564 $Y=-25360 $D=0
M924 BL<11> YOUT<3> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16379 $Y=-37036 $D=0
M925 BL<10> YOUT<2> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-16379 $Y=-27326 $D=0
M926 615 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-13645 $D=0
M927 BL<11> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-12110 $D=0
M928 616 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-10575 $D=0
M929 BL<11> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-9040 $D=0
M930 617 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-7505 $D=0
M931 BL<11> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-5970 $D=0
M932 618 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-4435 $D=0
M933 BL<11> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-2900 $D=0
M934 619 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=-1365 $D=0
M935 BL<11> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=170 $D=0
M936 620 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=1705 $D=0
M937 BL<11> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=3240 $D=0
M938 621 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=4775 $D=0
M939 BL<11> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=6310 $D=0
M940 622 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=7845 $D=0
M941 BL<11> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=9380 $D=0
M942 623 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=11335 $D=0
M943 BL<11> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=12870 $D=0
M944 624 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=14405 $D=0
M945 BL<11> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=15940 $D=0
M946 625 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=17475 $D=0
M947 BL<11> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=19010 $D=0
M948 626 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=20545 $D=0
M949 BL<11> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=22080 $D=0
M950 627 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=23615 $D=0
M951 BL<11> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=25150 $D=0
M952 628 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=26685 $D=0
M953 BL<11> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=28220 $D=0
M954 629 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=29755 $D=0
M955 BL<11> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=31290 $D=0
M956 630 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=32825 $D=0
M957 BL<11> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=34360 $D=0
M958 631 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=36315 $D=0
M959 BL<11> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=37850 $D=0
M960 632 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=39385 $D=0
M961 BL<11> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=40920 $D=0
M962 633 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=42455 $D=0
M963 BL<11> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=43990 $D=0
M964 634 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=45525 $D=0
M965 BL<11> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=47060 $D=0
M966 635 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=48595 $D=0
M967 BL<11> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=50130 $D=0
M968 636 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=51665 $D=0
M969 BL<11> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=53200 $D=0
M970 637 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=54735 $D=0
M971 BL<11> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=56270 $D=0
M972 638 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=57805 $D=0
M973 BL<11> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=59340 $D=0
M974 639 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=61295 $D=0
M975 BL<11> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=62830 $D=0
M976 640 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=64365 $D=0
M977 BL<11> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=65900 $D=0
M978 641 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=67435 $D=0
M979 BL<11> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=68970 $D=0
M980 642 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=70505 $D=0
M981 BL<11> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=72040 $D=0
M982 643 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=73575 $D=0
M983 BL<11> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=75110 $D=0
M984 644 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=76645 $D=0
M985 BL<11> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=78180 $D=0
M986 645 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=79715 $D=0
M987 BL<11> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=81250 $D=0
M988 646 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=82785 $D=0
M989 BL<11> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-16220 $Y=84320 $D=0
M990 VSS WL<63> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-13645 $D=0
M991 VSS WL<62> 647 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-12110 $D=0
M992 VSS WL<61> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-10575 $D=0
M993 VSS WL<60> 648 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-9040 $D=0
M994 VSS WL<59> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-7505 $D=0
M995 VSS WL<58> 649 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-5970 $D=0
M996 VSS WL<57> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-4435 $D=0
M997 VSS WL<56> 650 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-2900 $D=0
M998 VSS WL<55> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=-1365 $D=0
M999 VSS WL<54> 651 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=170 $D=0
M1000 VSS WL<53> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=1705 $D=0
M1001 VSS WL<52> 652 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=3240 $D=0
M1002 VSS WL<51> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=4775 $D=0
M1003 VSS WL<50> 653 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=6310 $D=0
M1004 VSS WL<49> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=7845 $D=0
M1005 VSS WL<48> 654 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=9380 $D=0
M1006 VSS WL<47> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=11335 $D=0
M1007 VSS WL<46> 655 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=12870 $D=0
M1008 VSS WL<45> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=14405 $D=0
M1009 VSS WL<44> 656 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=15940 $D=0
M1010 VSS WL<43> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=17475 $D=0
M1011 VSS WL<42> 657 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=19010 $D=0
M1012 VSS WL<41> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=20545 $D=0
M1013 VSS WL<40> 658 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=22080 $D=0
M1014 VSS WL<39> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=23615 $D=0
M1015 VSS WL<38> 659 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=25150 $D=0
M1016 VSS WL<37> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=26685 $D=0
M1017 VSS WL<36> 660 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=28220 $D=0
M1018 VSS WL<35> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=29755 $D=0
M1019 VSS WL<34> 661 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=31290 $D=0
M1020 VSS WL<33> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=32825 $D=0
M1021 VSS WL<32> 662 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=34360 $D=0
M1022 VSS WL<31> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=36315 $D=0
M1023 VSS WL<30> 663 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=37850 $D=0
M1024 VSS WL<29> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=39385 $D=0
M1025 VSS WL<28> 664 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=40920 $D=0
M1026 VSS WL<27> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=42455 $D=0
M1027 VSS WL<26> 665 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=43990 $D=0
M1028 VSS WL<25> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=45525 $D=0
M1029 VSS WL<24> 666 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=47060 $D=0
M1030 VSS WL<23> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=48595 $D=0
M1031 VSS WL<22> 667 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=50130 $D=0
M1032 VSS WL<21> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=51665 $D=0
M1033 VSS WL<20> 668 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=53200 $D=0
M1034 VSS WL<19> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=54735 $D=0
M1035 VSS WL<18> 669 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=56270 $D=0
M1036 VSS WL<17> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=57805 $D=0
M1037 VSS WL<16> 670 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=59340 $D=0
M1038 VSS WL<15> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=61295 $D=0
M1039 VSS WL<14> 671 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=62830 $D=0
M1040 VSS WL<13> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=64365 $D=0
M1041 VSS WL<12> 672 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=65900 $D=0
M1042 VSS WL<11> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=67435 $D=0
M1043 VSS WL<10> 673 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=68970 $D=0
M1044 VSS WL<9> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=70505 $D=0
M1045 VSS WL<8> 674 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=72040 $D=0
M1046 VSS WL<7> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=73575 $D=0
M1047 VSS WL<6> 675 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=75110 $D=0
M1048 VSS WL<5> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=76645 $D=0
M1049 VSS WL<4> 676 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=78180 $D=0
M1050 VSS WL<3> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=79715 $D=0
M1051 VSS WL<2> 677 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=81250 $D=0
M1052 VSS WL<1> BL<12> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=82785 $D=0
M1053 VSS WL<0> 678 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-14760 $Y=84320 $D=0
M1054 142 YOUT<5> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14414 $Y=-35070 $D=0
M1055 143 YOUT<4> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14414 $Y=-25360 $D=0
M1056 BL<13> YOUT<5> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14229 $Y=-37036 $D=0
M1057 BL<12> YOUT<4> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-14229 $Y=-27326 $D=0
M1058 679 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-13645 $D=0
M1059 BL<13> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-12110 $D=0
M1060 680 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-10575 $D=0
M1061 BL<13> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-9040 $D=0
M1062 681 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-7505 $D=0
M1063 BL<13> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-5970 $D=0
M1064 682 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-4435 $D=0
M1065 BL<13> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-2900 $D=0
M1066 683 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=-1365 $D=0
M1067 BL<13> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=170 $D=0
M1068 684 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=1705 $D=0
M1069 BL<13> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=3240 $D=0
M1070 685 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=4775 $D=0
M1071 BL<13> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=6310 $D=0
M1072 686 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=7845 $D=0
M1073 BL<13> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=9380 $D=0
M1074 687 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=11335 $D=0
M1075 BL<13> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=12870 $D=0
M1076 688 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=14405 $D=0
M1077 BL<13> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=15940 $D=0
M1078 689 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=17475 $D=0
M1079 BL<13> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=19010 $D=0
M1080 690 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=20545 $D=0
M1081 BL<13> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=22080 $D=0
M1082 691 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=23615 $D=0
M1083 BL<13> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=25150 $D=0
M1084 692 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=26685 $D=0
M1085 BL<13> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=28220 $D=0
M1086 693 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=29755 $D=0
M1087 BL<13> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=31290 $D=0
M1088 694 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=32825 $D=0
M1089 BL<13> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=34360 $D=0
M1090 695 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=36315 $D=0
M1091 BL<13> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=37850 $D=0
M1092 696 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=39385 $D=0
M1093 BL<13> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=40920 $D=0
M1094 697 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=42455 $D=0
M1095 BL<13> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=43990 $D=0
M1096 698 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=45525 $D=0
M1097 BL<13> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=47060 $D=0
M1098 699 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=48595 $D=0
M1099 BL<13> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=50130 $D=0
M1100 700 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=51665 $D=0
M1101 BL<13> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=53200 $D=0
M1102 701 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=54735 $D=0
M1103 BL<13> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=56270 $D=0
M1104 702 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=57805 $D=0
M1105 BL<13> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=59340 $D=0
M1106 703 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=61295 $D=0
M1107 BL<13> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=62830 $D=0
M1108 704 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=64365 $D=0
M1109 BL<13> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=65900 $D=0
M1110 705 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=67435 $D=0
M1111 BL<13> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=68970 $D=0
M1112 706 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=70505 $D=0
M1113 BL<13> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=72040 $D=0
M1114 707 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=73575 $D=0
M1115 BL<13> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=75110 $D=0
M1116 708 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=76645 $D=0
M1117 BL<13> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=78180 $D=0
M1118 709 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=79715 $D=0
M1119 BL<13> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=81250 $D=0
M1120 710 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=82785 $D=0
M1121 BL<13> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-14070 $Y=84320 $D=0
M1122 VSS WL<63> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-13645 $D=0
M1123 VSS WL<62> 711 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-12110 $D=0
M1124 VSS WL<61> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-10575 $D=0
M1125 VSS WL<60> 712 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-9040 $D=0
M1126 VSS WL<59> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-7505 $D=0
M1127 VSS WL<58> 713 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-5970 $D=0
M1128 VSS WL<57> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-4435 $D=0
M1129 VSS WL<56> 714 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-2900 $D=0
M1130 VSS WL<55> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=-1365 $D=0
M1131 VSS WL<54> 715 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=170 $D=0
M1132 VSS WL<53> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=1705 $D=0
M1133 VSS WL<52> 716 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=3240 $D=0
M1134 VSS WL<51> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=4775 $D=0
M1135 VSS WL<50> 717 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=6310 $D=0
M1136 VSS WL<49> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=7845 $D=0
M1137 VSS WL<48> 718 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=9380 $D=0
M1138 VSS WL<47> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=11335 $D=0
M1139 VSS WL<46> 719 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=12870 $D=0
M1140 VSS WL<45> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=14405 $D=0
M1141 VSS WL<44> 720 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=15940 $D=0
M1142 VSS WL<43> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=17475 $D=0
M1143 VSS WL<42> 721 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=19010 $D=0
M1144 VSS WL<41> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=20545 $D=0
M1145 VSS WL<40> 722 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=22080 $D=0
M1146 VSS WL<39> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=23615 $D=0
M1147 VSS WL<38> 723 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=25150 $D=0
M1148 VSS WL<37> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=26685 $D=0
M1149 VSS WL<36> 724 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=28220 $D=0
M1150 VSS WL<35> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=29755 $D=0
M1151 VSS WL<34> 725 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=31290 $D=0
M1152 VSS WL<33> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=32825 $D=0
M1153 VSS WL<32> 726 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=34360 $D=0
M1154 VSS WL<31> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=36315 $D=0
M1155 VSS WL<30> 727 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=37850 $D=0
M1156 VSS WL<29> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=39385 $D=0
M1157 VSS WL<28> 728 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=40920 $D=0
M1158 VSS WL<27> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=42455 $D=0
M1159 VSS WL<26> 729 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=43990 $D=0
M1160 VSS WL<25> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=45525 $D=0
M1161 VSS WL<24> 730 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=47060 $D=0
M1162 VSS WL<23> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=48595 $D=0
M1163 VSS WL<22> 731 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=50130 $D=0
M1164 VSS WL<21> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=51665 $D=0
M1165 VSS WL<20> 732 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=53200 $D=0
M1166 VSS WL<19> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=54735 $D=0
M1167 VSS WL<18> 733 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=56270 $D=0
M1168 VSS WL<17> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=57805 $D=0
M1169 VSS WL<16> 734 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=59340 $D=0
M1170 VSS WL<15> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=61295 $D=0
M1171 VSS WL<14> 735 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=62830 $D=0
M1172 VSS WL<13> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=64365 $D=0
M1173 VSS WL<12> 736 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=65900 $D=0
M1174 VSS WL<11> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=67435 $D=0
M1175 VSS WL<10> 737 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=68970 $D=0
M1176 VSS WL<9> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=70505 $D=0
M1177 VSS WL<8> 738 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=72040 $D=0
M1178 VSS WL<7> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=73575 $D=0
M1179 VSS WL<6> 739 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=75110 $D=0
M1180 VSS WL<5> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=76645 $D=0
M1181 VSS WL<4> 740 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=78180 $D=0
M1182 VSS WL<3> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=79715 $D=0
M1183 VSS WL<2> 741 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=81250 $D=0
M1184 VSS WL<1> BL<14> VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=82785 $D=0
M1185 VSS WL<0> 742 VSS N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06 $X=-12610 $Y=84320 $D=0
M1186 144 YOUT<7> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12264 $Y=-35070 $D=0
M1187 145 YOUT<6> VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12264 $Y=-25360 $D=0
M1188 BL<15> YOUT<7> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12079 $Y=-37036 $D=0
M1189 BL<14> YOUT<6> DL<1> VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-12079 $Y=-27326 $D=0
M1190 743 WL<63> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-13645 $D=0
M1191 BL<15> WL<62> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-12110 $D=0
M1192 744 WL<61> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-10575 $D=0
M1193 BL<15> WL<60> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-9040 $D=0
M1194 745 WL<59> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-7505 $D=0
M1195 BL<15> WL<58> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-5970 $D=0
M1196 746 WL<57> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-4435 $D=0
M1197 BL<15> WL<56> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-2900 $D=0
M1198 747 WL<55> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=-1365 $D=0
M1199 BL<15> WL<54> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=170 $D=0
M1200 748 WL<53> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=1705 $D=0
M1201 BL<15> WL<52> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=3240 $D=0
M1202 749 WL<51> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=4775 $D=0
M1203 BL<15> WL<50> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=6310 $D=0
M1204 750 WL<49> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=7845 $D=0
M1205 BL<15> WL<48> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=9380 $D=0
M1206 751 WL<47> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=11335 $D=0
M1207 BL<15> WL<46> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=12870 $D=0
M1208 752 WL<45> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=14405 $D=0
M1209 BL<15> WL<44> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=15940 $D=0
M1210 753 WL<43> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=17475 $D=0
M1211 BL<15> WL<42> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=19010 $D=0
M1212 754 WL<41> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=20545 $D=0
M1213 BL<15> WL<40> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=22080 $D=0
M1214 755 WL<39> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=23615 $D=0
M1215 BL<15> WL<38> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=25150 $D=0
M1216 756 WL<37> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=26685 $D=0
M1217 BL<15> WL<36> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=28220 $D=0
M1218 757 WL<35> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=29755 $D=0
M1219 BL<15> WL<34> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=31290 $D=0
M1220 758 WL<33> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=32825 $D=0
M1221 BL<15> WL<32> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=34360 $D=0
M1222 759 WL<31> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=36315 $D=0
M1223 BL<15> WL<30> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=37850 $D=0
M1224 760 WL<29> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=39385 $D=0
M1225 BL<15> WL<28> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=40920 $D=0
M1226 761 WL<27> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=42455 $D=0
M1227 BL<15> WL<26> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=43990 $D=0
M1228 762 WL<25> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=45525 $D=0
M1229 BL<15> WL<24> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=47060 $D=0
M1230 763 WL<23> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=48595 $D=0
M1231 BL<15> WL<22> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=50130 $D=0
M1232 764 WL<21> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=51665 $D=0
M1233 BL<15> WL<20> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=53200 $D=0
M1234 765 WL<19> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=54735 $D=0
M1235 BL<15> WL<18> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=56270 $D=0
M1236 766 WL<17> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=57805 $D=0
M1237 BL<15> WL<16> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=59340 $D=0
M1238 767 WL<15> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=61295 $D=0
M1239 BL<15> WL<14> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=62830 $D=0
M1240 768 WL<13> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=64365 $D=0
M1241 BL<15> WL<12> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=65900 $D=0
M1242 769 WL<11> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=67435 $D=0
M1243 BL<15> WL<10> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=68970 $D=0
M1244 770 WL<9> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=70505 $D=0
M1245 BL<15> WL<8> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=72040 $D=0
M1246 771 WL<7> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=73575 $D=0
M1247 BL<15> WL<6> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=75110 $D=0
M1248 772 WL<5> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=76645 $D=0
M1249 BL<15> WL<4> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=78180 $D=0
M1250 773 WL<3> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=79715 $D=0
M1251 BL<15> WL<2> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=81250 $D=0
M1252 774 WL<1> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=82785 $D=0
M1253 BL<15> WL<0> VSS VSS N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07 $X=-11920 $Y=84320 $D=0
M1254 61 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=8965 $D=1
M1255 59 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=21005 $D=1
M1256 63 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=33045 $D=1
M1257 62 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=57645 $D=1
M1258 60 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=69685 $D=1
M1259 64 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-66670 $Y=81725 $D=1
M1260 16 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-11510 $D=1
M1261 16 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-10050 $D=1
M1262 16 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-8590 $D=1
M1263 16 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-7130 $D=1
M1264 17 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-5490 $D=1
M1265 17 61 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-4030 $D=1
M1266 17 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-2570 $D=1
M1267 17 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=-1110 $D=1
M1268 18 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=530 $D=1
M1269 18 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=1990 $D=1
M1270 18 59 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=3450 $D=1
M1271 18 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=4910 $D=1
M1272 19 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=6550 $D=1
M1273 19 61 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=8010 $D=1
M1274 19 59 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=9470 $D=1
M1275 19 X_sel<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=10930 $D=1
M1276 20 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=12570 $D=1
M1277 20 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=14030 $D=1
M1278 20 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=15490 $D=1
M1279 20 63 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=16950 $D=1
M1280 21 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=18590 $D=1
M1281 21 61 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=20050 $D=1
M1282 21 X_sel<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=21510 $D=1
M1283 21 63 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=22970 $D=1
M1284 22 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=24610 $D=1
M1285 22 X_sel<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=26070 $D=1
M1286 22 59 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=27530 $D=1
M1287 22 63 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=28990 $D=1
M1288 23 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=30630 $D=1
M1289 23 61 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=32090 $D=1
M1290 23 59 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=33550 $D=1
M1291 23 63 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=35010 $D=1
M1292 24 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=37170 $D=1
M1293 24 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=38630 $D=1
M1294 24 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=40090 $D=1
M1295 24 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=41550 $D=1
M1296 25 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=43190 $D=1
M1297 25 62 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=44650 $D=1
M1298 25 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=46110 $D=1
M1299 25 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=47570 $D=1
M1300 26 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=49210 $D=1
M1301 26 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=50670 $D=1
M1302 26 60 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=52130 $D=1
M1303 26 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=53590 $D=1
M1304 27 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=55230 $D=1
M1305 27 62 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=56690 $D=1
M1306 27 60 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=58150 $D=1
M1307 27 X_sel<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=59610 $D=1
M1308 28 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=61250 $D=1
M1309 28 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=62710 $D=1
M1310 28 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=64170 $D=1
M1311 28 64 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=65630 $D=1
M1312 29 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=67270 $D=1
M1313 29 62 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=68730 $D=1
M1314 29 X_sel<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=70190 $D=1
M1315 29 64 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=71650 $D=1
M1316 30 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=73290 $D=1
M1317 30 X_sel<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=74750 $D=1
M1318 30 60 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=76210 $D=1
M1319 30 64 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=77670 $D=1
M1320 31 WL_EN VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=79310 $D=1
M1321 31 62 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=80770 $D=1
M1322 31 60 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=82230 $D=1
M1323 31 64 VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-56945 $Y=83690 $D=1
M1324 WL<63> 16 199 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-13505 $D=1
M1325 WL<62> 16 200 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-11970 $D=1
M1326 WL<61> 16 201 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-10435 $D=1
M1327 WL<60> 16 202 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-8900 $D=1
M1328 WL<59> 16 203 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-7365 $D=1
M1329 WL<58> 16 204 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-5830 $D=1
M1330 WL<57> 16 205 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-4295 $D=1
M1331 WL<56> 16 206 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-2760 $D=1
M1332 WL<55> 17 207 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=-1225 $D=1
M1333 WL<54> 17 208 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=310 $D=1
M1334 WL<53> 17 209 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=1845 $D=1
M1335 WL<52> 17 210 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=3380 $D=1
M1336 WL<51> 17 211 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=4915 $D=1
M1337 WL<50> 17 212 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=6450 $D=1
M1338 WL<49> 17 213 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=7985 $D=1
M1339 WL<48> 17 214 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=9520 $D=1
M1340 WL<47> 18 215 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=11475 $D=1
M1341 WL<46> 18 216 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=13010 $D=1
M1342 WL<45> 18 217 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=14545 $D=1
M1343 WL<44> 18 218 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=16080 $D=1
M1344 WL<43> 18 219 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=17615 $D=1
M1345 WL<42> 18 220 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=19150 $D=1
M1346 WL<41> 18 221 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=20685 $D=1
M1347 WL<40> 18 222 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=22220 $D=1
M1348 WL<39> 19 223 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=23755 $D=1
M1349 WL<38> 19 224 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=25290 $D=1
M1350 WL<37> 19 225 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=26825 $D=1
M1351 WL<36> 19 226 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=28360 $D=1
M1352 WL<35> 19 227 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=29895 $D=1
M1353 WL<34> 19 228 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=31430 $D=1
M1354 WL<33> 19 229 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=32965 $D=1
M1355 WL<32> 19 230 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=34500 $D=1
M1356 WL<31> 20 231 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=36455 $D=1
M1357 WL<30> 20 232 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=37990 $D=1
M1358 WL<29> 20 233 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=39525 $D=1
M1359 WL<28> 20 234 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=41060 $D=1
M1360 WL<27> 20 235 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=42595 $D=1
M1361 WL<26> 20 236 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=44130 $D=1
M1362 WL<25> 20 237 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=45665 $D=1
M1363 WL<24> 20 238 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=47200 $D=1
M1364 WL<23> 21 239 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=48735 $D=1
M1365 WL<22> 21 240 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=50270 $D=1
M1366 WL<21> 21 241 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=51805 $D=1
M1367 WL<20> 21 242 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=53340 $D=1
M1368 WL<19> 21 243 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=54875 $D=1
M1369 WL<18> 21 244 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=56410 $D=1
M1370 WL<17> 21 245 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=57945 $D=1
M1371 WL<16> 21 246 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=59480 $D=1
M1372 WL<15> 22 247 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=61435 $D=1
M1373 WL<14> 22 248 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=62970 $D=1
M1374 WL<13> 22 249 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=64505 $D=1
M1375 WL<12> 22 250 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=66040 $D=1
M1376 WL<11> 22 251 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=67575 $D=1
M1377 WL<10> 22 252 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=69110 $D=1
M1378 WL<9> 22 253 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=70645 $D=1
M1379 WL<8> 22 254 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=72180 $D=1
M1380 WL<7> 23 255 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=73715 $D=1
M1381 WL<6> 23 256 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=75250 $D=1
M1382 WL<5> 23 257 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=76785 $D=1
M1383 WL<4> 23 258 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=78320 $D=1
M1384 WL<3> 23 259 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=79855 $D=1
M1385 WL<2> 23 260 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=81390 $D=1
M1386 WL<1> 23 261 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=82925 $D=1
M1387 WL<0> 23 262 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-37950 $Y=84460 $D=1
M1388 VDD 24 199 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-13505 $D=1
M1389 VDD 25 200 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-11970 $D=1
M1390 VDD 26 201 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-10435 $D=1
M1391 VDD 27 202 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-8900 $D=1
M1392 VDD 28 203 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-7365 $D=1
M1393 VDD 29 204 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-5830 $D=1
M1394 VDD 30 205 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-4295 $D=1
M1395 VDD 31 206 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-2760 $D=1
M1396 VDD 24 207 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=-1225 $D=1
M1397 VDD 25 208 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=310 $D=1
M1398 VDD 26 209 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=1845 $D=1
M1399 VDD 27 210 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=3380 $D=1
M1400 VDD 28 211 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=4915 $D=1
M1401 VDD 29 212 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=6450 $D=1
M1402 VDD 30 213 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=7985 $D=1
M1403 VDD 31 214 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=9520 $D=1
M1404 VDD 24 215 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=11475 $D=1
M1405 VDD 25 216 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=13010 $D=1
M1406 VDD 26 217 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=14545 $D=1
M1407 VDD 27 218 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=16080 $D=1
M1408 VDD 28 219 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=17615 $D=1
M1409 VDD 29 220 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=19150 $D=1
M1410 VDD 30 221 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=20685 $D=1
M1411 VDD 31 222 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=22220 $D=1
M1412 VDD 24 223 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=23755 $D=1
M1413 VDD 25 224 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=25290 $D=1
M1414 VDD 26 225 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=26825 $D=1
M1415 VDD 27 226 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=28360 $D=1
M1416 VDD 28 227 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=29895 $D=1
M1417 VDD 29 228 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=31430 $D=1
M1418 VDD 30 229 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=32965 $D=1
M1419 VDD 31 230 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=34500 $D=1
M1420 VDD 24 231 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=36455 $D=1
M1421 VDD 25 232 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=37990 $D=1
M1422 VDD 26 233 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=39525 $D=1
M1423 VDD 27 234 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=41060 $D=1
M1424 VDD 28 235 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=42595 $D=1
M1425 VDD 29 236 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=44130 $D=1
M1426 VDD 30 237 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=45665 $D=1
M1427 VDD 31 238 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=47200 $D=1
M1428 VDD 24 239 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=48735 $D=1
M1429 VDD 25 240 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=50270 $D=1
M1430 VDD 26 241 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=51805 $D=1
M1431 VDD 27 242 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=53340 $D=1
M1432 VDD 28 243 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=54875 $D=1
M1433 VDD 29 244 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=56410 $D=1
M1434 VDD 30 245 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=57945 $D=1
M1435 VDD 31 246 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=59480 $D=1
M1436 VDD 24 247 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=61435 $D=1
M1437 VDD 25 248 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=62970 $D=1
M1438 VDD 26 249 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=64505 $D=1
M1439 VDD 27 250 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=66040 $D=1
M1440 VDD 28 251 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=67575 $D=1
M1441 VDD 29 252 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=69110 $D=1
M1442 VDD 30 253 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=70645 $D=1
M1443 VDD 31 254 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=72180 $D=1
M1444 VDD 24 255 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=73715 $D=1
M1445 VDD 25 256 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=75250 $D=1
M1446 VDD 26 257 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=76785 $D=1
M1447 VDD 27 258 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=78320 $D=1
M1448 VDD 28 259 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=79855 $D=1
M1449 VDD 29 260 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=81390 $D=1
M1450 VDD 30 261 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=82925 $D=1
M1451 VDD 31 262 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=-35145 $Y=84460 $D=1
M1452 VDD CLK BL<0> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-27660 $Y=-17045 $D=1
M1453 130 YOUT<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-33365 $D=1
M1454 DL<0> 130 BL<1> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-30465 $D=1
M1455 131 YOUT<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-23655 $D=1
M1456 DL<0> 131 BL<0> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-27314 $Y=-20755 $D=1
M1457 BL<1> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-26970 $Y=-17045 $D=1
M1458 VDD CLK BL<2> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-25510 $Y=-17045 $D=1
M1459 132 YOUT<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-25164 $Y=-33365 $D=1
M1460 DL<0> 132 BL<3> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-25164 $Y=-30465 $D=1
M1461 133 YOUT<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-25164 $Y=-23655 $D=1
M1462 DL<0> 133 BL<2> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-25164 $Y=-20755 $D=1
M1463 BL<3> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-24820 $Y=-17045 $D=1
M1464 VDD CLK BL<4> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-23360 $Y=-17045 $D=1
M1465 134 YOUT<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-33365 $D=1
M1466 DL<0> 134 BL<5> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-30465 $D=1
M1467 135 YOUT<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-23655 $D=1
M1468 DL<0> 135 BL<4> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-23014 $Y=-20755 $D=1
M1469 BL<5> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-22670 $Y=-17045 $D=1
M1470 VDD CLK BL<6> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-21210 $Y=-17045 $D=1
M1471 136 YOUT<7> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-33365 $D=1
M1472 DL<0> 136 BL<7> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-30465 $D=1
M1473 137 YOUT<6> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-23655 $D=1
M1474 DL<0> 137 BL<6> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-20864 $Y=-20755 $D=1
M1475 BL<7> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-20520 $Y=-17045 $D=1
M1476 VDD CLK BL<8> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-19060 $Y=-17045 $D=1
M1477 138 YOUT<1> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-33365 $D=1
M1478 DL<1> 138 BL<9> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-30465 $D=1
M1479 139 YOUT<0> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-23655 $D=1
M1480 DL<1> 139 BL<8> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-18714 $Y=-20755 $D=1
M1481 BL<9> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-18370 $Y=-17045 $D=1
M1482 VDD CLK BL<10> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-16910 $Y=-17045 $D=1
M1483 140 YOUT<3> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-33365 $D=1
M1484 DL<1> 140 BL<11> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-30465 $D=1
M1485 141 YOUT<2> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-23655 $D=1
M1486 DL<1> 141 BL<10> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-16564 $Y=-20755 $D=1
M1487 BL<11> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-16220 $Y=-17045 $D=1
M1488 VDD CLK BL<12> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-14760 $Y=-17045 $D=1
M1489 142 YOUT<5> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-33365 $D=1
M1490 DL<1> 142 BL<13> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-30465 $D=1
M1491 143 YOUT<4> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-23655 $D=1
M1492 DL<1> 143 BL<12> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-14414 $Y=-20755 $D=1
M1493 BL<13> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-14070 $Y=-17045 $D=1
M1494 VDD CLK BL<14> VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=-12610 $Y=-17045 $D=1
M1495 144 YOUT<7> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-33365 $D=1
M1496 DL<1> 144 BL<15> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-30465 $D=1
M1497 145 YOUT<6> VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-23655 $D=1
M1498 DL<1> 145 BL<14> VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-12264 $Y=-20755 $D=1
M1499 BL<15> CLK VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=-11920 $Y=-17045 $D=1
X1500 Dout<0> SO<0> SAEN DL<0> VSS Vref VDD Final_SA $T=-23415 -43080 0 0 $X=-26580 $Y=-45535
X1501 Dout<1> SO<1> SAEN DL<1> VSS Vref VDD Final_SA $T=-15255 -43080 0 0 $X=-18420 $Y=-45535
X1502 CLK VSS VDD 9 inv_final $T=-68030 -26395 0 0 $X=-69190 $Y=-29660
X1503 776 VSS VDD 148 inv_final $T=-65830 -33650 0 0 $X=-66990 $Y=-36915
X1504 CLK 146 VDD VSS WL_EN final_and $T=-54685 -45770 0 0 $X=-47930 $Y=-46920
X1505 CLK 65 VDD VSS SAEN final_and $T=-44075 -45770 0 0 $X=-37320 $Y=-46920
X1506 777 VSS VDD 778 776 ICV_1 $T=-69030 -33650 0 0 $X=-70190 $Y=-36915
X1507 148 VSS VDD 779 780 ICV_2 $T=-88270 -43555 0 0 $X=-89430 $Y=-46820
X1508 CLK VSS VDD 781 782 ICV_2 $T=-88230 -33650 0 0 $X=-89390 $Y=-36915
X1509 780 VSS VDD 783 784 ICV_2 $T=-81870 -43555 0 0 $X=-83030 $Y=-46820
X1510 782 VSS VDD 785 786 ICV_2 $T=-81830 -33650 0 0 $X=-82990 $Y=-36915
X1511 784 VSS VDD 787 788 ICV_2 $T=-75470 -43555 0 0 $X=-76630 $Y=-46820
X1512 786 VSS VDD 789 777 ICV_2 $T=-75430 -33650 0 0 $X=-76590 $Y=-36915
X1513 788 VSS VDD 790 791 ICV_2 $T=-69070 -43555 0 0 $X=-70230 $Y=-46820
X1514 791 VSS VDD 792 793 ICV_2 $T=-62670 -43555 0 0 $X=-63830 $Y=-46820
X1515 793 VSS VDD 65 146 ICV_2 $T=-56270 -43555 0 0 $X=-57430 $Y=-46820
X1516 Y_sel<0> Y_sel<1> Y_sel<2> YOUT<3> YOUT<2> YOUT<1> YOUT<0> YOUT<7> YOUT<6> YOUT<5> YOUT<4> VDD VSS Ydecoder_final $T=-62420 -36975 0 0 $X=-62800 $Y=-40160
X1517 9 CLK VSS VDD A<2> Y_sel<2> FInal_FF $T=-84440 -21020 0 0 $X=-90065 $Y=-28235
X1518 9 CLK VSS VDD A<1> Y_sel<1> FInal_FF $T=-84440 -8310 0 0 $X=-90065 $Y=-15525
X1519 9 CLK VSS VDD A<0> Y_sel<0> FInal_FF $T=-84440 4400 0 0 $X=-90065 $Y=-2815
X1520 9 CLK VSS VDD A<6> X_sel<3> FInal_FF $T=-84440 17110 0 0 $X=-90065 $Y=9895
X1521 9 CLK VSS VDD A<7> X_sel<4> FInal_FF $T=-84440 29820 0 0 $X=-90065 $Y=22605
X1522 9 CLK VSS VDD A<8> X_sel<5> FInal_FF $T=-84440 42530 0 0 $X=-90065 $Y=35315
X1523 9 CLK VSS VDD A<3> X_sel<0> FInal_FF $T=-84440 55240 0 0 $X=-90065 $Y=48025
X1524 9 CLK VSS VDD A<4> X_sel<1> FInal_FF $T=-84440 67950 0 0 $X=-90065 $Y=60735
X1525 9 CLK VSS VDD A<5> X_sel<2> FInal_FF $T=-84440 80660 0 0 $X=-90065 $Y=73445
.ENDS
***************************************
