************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: hw2_part1_1
* View Name:     schematic
* Netlisted on:  Nov  5 08:47:54 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    hw2_part1_1
* View Name:    schematic
************************************************************************

.SUBCKT hw2_part1_1 A B C OUT VDD VSS
*.PININFO A:I B:I C:I OUT:O VDD:B VSS:B
MM6 net6 C VSS VSS N_18 W=2u L=180.00n m=4
MM5 net10 B net6 VSS N_18 W=2u L=180.00n m=4
MM4 OUT A net10 VSS N_18 W=2u L=180.00n m=4
MM2 OUT C VDD VDD P_18 W=1.5u L=180.00n m=1
MM1 OUT A VDD VDD P_18 W=1.5u L=180.00n m=10
MM0 OUT B VDD VDD P_18 W=1.5u L=180.00n m=1
.ENDS

