* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT inv_1u5_0u5 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 4 1 2 2 N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-65 $Y=-2195 $D=0
M1 4 1 3 3 P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-65 $Y=-490 $D=1
.ENDS
***************************************
.SUBCKT FInal_FF !c C VSS VDD D Q
** N=15 EP=6 IP=16 FDC=20
M0 7 !c 4 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=-2285 $Y=-2400 $D=0
M1 9 C VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=1670 $Y=-2400 $D=0
M2 4 10 9 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=3170 $Y=-2400 $D=0
M3 5 C 10 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=5540 $Y=-1425 $D=0
M4 11 !c VSS VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=9425 $Y=-2400 $D=0
M5 5 13 11 VSS N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=2.55e-13 PD=1.52e-06 PS=1.52e-06 $X=10925 $Y=-2400 $D=0
M6 7 C 4 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=-2285 $Y=-5120 $D=1
M7 8 !c VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=1570 $Y=-5120 $D=1
M8 4 10 8 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=3170 $Y=-5120 $D=1
M9 5 !c 10 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=5540 $Y=295 $D=1
M10 12 C VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=9425 $Y=-5120 $D=1
M11 5 13 12 VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=7.65e-13 PD=2.52e-06 PS=2.52e-06 $X=10925 $Y=-5120 $D=1
X12 D VSS VDD 7 inv_1u5_0u5 $T=-2220 1570 0 0 $X=-3380 $Y=-1695
X13 4 VSS VDD 10 inv_1u5_0u5 $T=1735 1565 0 0 $X=575 $Y=-1700
X14 5 VSS VDD 13 inv_1u5_0u5 $T=9490 1565 0 0 $X=8330 $Y=-1700
X15 13 VSS VDD Q inv_1u5_0u5 $T=13725 1565 0 0 $X=12565 $Y=-1700
.ENDS
***************************************
