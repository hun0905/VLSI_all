************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: 3to8decoder_en
* View Name:     schematic
* Netlisted on:  Jan 12 17:52:21 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    nand4
* View Name:    schematic
************************************************************************

.SUBCKT nand4 A B C D OUT VDD VSS
*.PININFO A:I B:I C:I D:I OUT:O VDD:B VSS:B
MM11 net030 D VSS VSS N_18 W=500.0n L=180.00n m=1
MM6 net40 C net030 VSS N_18 W=500.0n L=180.00n m=1
MM5 net44 B net40 VSS N_18 W=500.0n L=180.00n m=1
MM4 OUT A net44 VSS N_18 W=500.0n L=180.00n m=1
MM12 OUT D VDD VDD P_18 W=500.0n L=180.00n m=3
MM10 OUT A VDD VDD P_18 W=500.0n L=180.00n m=3
MM2 OUT C VDD VDD P_18 W=500.0n L=180.00n m=3
MM0 OUT B VDD VDD P_18 W=500.0n L=180.00n m=3
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter IN OUT VDD VSS
*.PININFO IN:I OUT:B VDD:B VSS:B
MM10 OUT IN VSS VSS N_18 W=500.0n L=180.00n m=1
MM6 OUT IN VDD VDD P_18 W=1.5u L=180.00n m=1
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    3to8decoder_en
* View Name:    schematic
************************************************************************

.SUBCKT 3to8decoder_en A B C EN OUT0 OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 OUT7 VDD VSS
*.PININFO A:I B:I C:I EN:I OUT0:O OUT1:O OUT2:O OUT3:O OUT4:O OUT5:O OUT6:O 
*.PININFO OUT7:O VDD:B VSS:B
XI7 A B C EN OUT7 VDD VSS / nand4
XI6 A B net0116 EN OUT6 VDD VSS / nand4
XI5 A net0105 C EN OUT5 VDD VSS / nand4
XI4 A net0105 net0116 EN OUT4 VDD VSS / nand4
XI3 net0158 B C EN OUT3 VDD VSS / nand4
XI2 net0158 B net0116 EN OUT2 VDD VSS / nand4
XI1 net0158 net0105 C EN OUT1 VDD VSS / nand4
XI0 net0158 net0105 net0116 EN OUT0 VDD VSS / nand4
XI11 B net0105 VDD VSS / inverter
XI10 C net0116 VDD VSS / inverter
XI8 A net0158 VDD VSS / inverter
.ENDS

