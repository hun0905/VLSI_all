************************************************************************
* auCdl Netlist:
* 
* Library Name:  vlsi
* Top Cell Name: Final_noSA
* View Name:     schematic
* Netlisted on:  Jan 16 20:32:49 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: vlsi
* Cell Name:    and
* View Name:    schematic
************************************************************************

.SUBCKT and A B OUT VDD VSS
*.PININFO A:I B:I OUT:O VDD:B VSS:B
MM10 OUT net067 VSS VSS N_18 W=500.0n L=180.00n m=1
MM5 net44 B VSS VSS N_18 W=500.0n L=180.00n m=1
MM4 net067 A net44 VSS N_18 W=500.0n L=180.00n m=1
MM9 OUT net067 VDD VDD P_18 W=500.0n L=180.00n m=3
MM1 net067 A VDD VDD P_18 W=500.0n L=180.00n m=3
MM0 net067 B VDD VDD P_18 W=500.0n L=180.00n m=3
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter IN OUT VDD VSS
*.PININFO IN:I OUT:B VDD:B VSS:B
MM10 OUT IN VSS VSS N_18 W=500.0n L=180.00n m=1
MM6 OUT IN VDD VDD P_18 W=1.5u L=180.00n m=1
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    buffer
* View Name:    schematic
************************************************************************

.SUBCKT buffer IN OUT VDD VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
XI7 net14 OUT VDD VSS / inverter
XI5 IN net14 VDD VSS / inverter
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    tri_state
* View Name:    schematic
************************************************************************

.SUBCKT tri_state !en VDD VSS en input out
*.PININFO !en:I VDD:I VSS:I en:I input:I out:B
MM3 net5 en VSS VSS N_18 W=500.0n L=180.00n
MM2 out input net5 VSS N_18 W=500.0n L=180.00n
MM1 out input net12 VDD P_18 W=1.5u L=180.00n
MM0 net12 !en VDD VDD P_18 W=1.5u L=180.00n
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    Final_FF
* View Name:    schematic
************************************************************************

.SUBCKT Final_FF !c C D Q VDD VSS
*.PININFO !c:I C:I D:I Q:O VDD:B VSS:B
MM4 net5 C net14 VSS N_18 W=500.0n L=180.00n
MM2 net18 !c net13 VSS N_18 W=500.0n L=180.00n
MM3 net5 !c net14 VDD P_18 W=1.5u L=180.00n
MM0 net18 C net13 VDD P_18 W=1.5u L=180.00n
XI6 C VDD VSS !c net1 net5 / tri_state
XI5 !c VDD VSS C net14 net13 / tri_state
XI4 net1 Q VDD VSS / inverter
XI3 net5 net1 VDD VSS / inverter
XI1 net13 net14 VDD VSS / inverter
XI0 D net18 VDD VSS / inverter
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    timing_control2
* View Name:    schematic
************************************************************************

.SUBCKT timing_control2 A<0> A<1> A<2> A<3> A<4> A<5> A<6> A<7> A<8> CLK SAEN 
+ VDD VSS WL_EN X_sel_FF<0> X_sel_FF<1> X_sel_FF<2> X_sel_FF<3> X_sel_FF<4> 
+ X_sel_FF<5> Y_sel_FF<0> Y_sel_FF<1> Y_sel_FF<2>
*.PININFO A<0>:I A<1>:I A<2>:I A<3>:I A<4>:I A<5>:I A<6>:I A<7>:I A<8>:I CLK:I 
*.PININFO SAEN:O WL_EN:O X_sel_FF<0>:O X_sel_FF<1>:O X_sel_FF<2>:O 
*.PININFO X_sel_FF<3>:O X_sel_FF<4>:O X_sel_FF<5>:O Y_sel_FF<0>:O 
*.PININFO Y_sel_FF<1>:O Y_sel_FF<2>:O VDD:B VSS:B
XI43 CLK net0134 SAEN VDD VSS / and
XI42 CLK net101 WL_EN VDD VSS / and
XI60 net0134 net101 VDD VSS / inverter
XI44 CLK net0145 VDD VSS / inverter
XI61 net0170 net092 VDD VSS / buffer
XI63 net092 net099 VDD VSS / buffer
XI65 net099 net0134 VDD VSS / buffer
XI69 net097 net096 VDD VSS / buffer
XI70 net0182 net097 VDD VSS / buffer
XI71 net0162 net0158 VDD VSS / buffer
XI72 net0185 net0162 VDD VSS / buffer
XI74 net0174 net0170 VDD VSS / buffer
XI75 net096 net0174 VDD VSS / buffer
XI77 net0158 net0182 VDD VSS / buffer
XI50 net0146 net094 VDD VSS / buffer
XI55 net0142 net098 VDD VSS / buffer
XI51 net094 net0102 VDD VSS / buffer
XI58 net0114 net0106 VDD VSS / buffer
XI52 net0102 net0110 VDD VSS / buffer
XI57 net0118 net0114 VDD VSS / buffer
XI56 net098 net0118 VDD VSS / buffer
XI59 net0106 net0185 VDD VSS / buffer
XI47 net0130 net0126 VDD VSS / buffer
XI46 net113 net0130 VDD VSS / buffer
XI39 net109 net105 VDD VSS / buffer
XI38 CLK net109 VDD VSS / buffer
XI54 net0154 net0142 VDD VSS / buffer
XI49 net0150 net0146 VDD VSS / buffer
XI48 net0126 net0150 VDD VSS / buffer
XI53 net0110 net0154 VDD VSS / buffer
XI40 net105 net113 VDD VSS / buffer
XI21 net0145 CLK A<8> X_sel_FF<5> VDD VSS / Final_FF
XI29 net0145 CLK A<5> X_sel_FF<2> VDD VSS / Final_FF
XI28 net0145 CLK A<7> X_sel_FF<4> VDD VSS / Final_FF
XI30 net0145 CLK A<6> X_sel_FF<3> VDD VSS / Final_FF
XI31 net0145 CLK A<2> Y_sel_FF<2> VDD VSS / Final_FF
XI32 net0145 CLK A<1> Y_sel_FF<1> VDD VSS / Final_FF
XI33 net0145 CLK A<3> X_sel_FF<0> VDD VSS / Final_FF
XI34 net0145 CLK A<4> X_sel_FF<1> VDD VSS / Final_FF
XI35 net0145 CLK A<0> Y_sel_FF<0> VDD VSS / Final_FF
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    SA_Final
* View Name:    schematic
************************************************************************

.SUBCKT SA_Final EN INN INP SO SON VDD VSS
*.PININFO EN:I INN:I INP:I SO:O SON:O VDD:B VSS:B
MM19 net096 EN VSS VSS N_18 W=500.0n L=180.00n m=4
MM17 SON SO net089 VSS N_18 W=500.0n L=180.00n m=1
MM18 net089 INP net096 VSS N_18 W=500.0n L=180.00n m=1
MM16 net093 INN net096 VSS N_18 W=500.0n L=180.00n m=1
MM15 SO SON net093 VSS N_18 W=500.0n L=180.00n m=1
MM13 SON SO VDD VDD P_18 W=500.0n L=180.00n m=1
MM12 SO SON VDD VDD P_18 W=500.0n L=180.00n m=1
MM9 SON EN VDD VDD P_18 W=500.0n L=180.00n m=1
MM11 SO EN VDD VDD P_18 W=500.0n L=180.00n m=1
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    nand4
* View Name:    schematic
************************************************************************

.SUBCKT nand4 A B C D OUT VDD VSS
*.PININFO A:I B:I C:I D:I OUT:O VDD:B VSS:B
MM11 net030 D VSS VSS N_18 W=500.0n L=180.00n m=1
MM6 net40 C net030 VSS N_18 W=500.0n L=180.00n m=1
MM5 net44 B net40 VSS N_18 W=500.0n L=180.00n m=1
MM4 OUT A net44 VSS N_18 W=500.0n L=180.00n m=1
MM12 OUT D VDD VDD P_18 W=500.0n L=180.00n m=3
MM10 OUT A VDD VDD P_18 W=500.0n L=180.00n m=3
MM2 OUT C VDD VDD P_18 W=500.0n L=180.00n m=3
MM0 OUT B VDD VDD P_18 W=500.0n L=180.00n m=3
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    3to8decoder_en
* View Name:    schematic
************************************************************************

.SUBCKT to8decoder_en A B C EN OUT0 OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 OUT7 VDD VSS
*.PININFO A:I B:I C:I EN:I OUT0:O OUT1:O OUT2:O OUT3:O OUT4:O OUT5:O OUT6:O 
*.PININFO OUT7:O VDD:B VSS:B
XI7 A B C EN OUT7 VDD VSS / nand4
XI6 A B net0116 EN OUT6 VDD VSS / nand4
XI5 A net0105 C EN OUT5 VDD VSS / nand4
XI4 A net0105 net0116 EN OUT4 VDD VSS / nand4
XI3 net0158 B C EN OUT3 VDD VSS / nand4
XI2 net0158 B net0116 EN OUT2 VDD VSS / nand4
XI1 net0158 net0105 C EN OUT1 VDD VSS / nand4
XI0 net0158 net0105 net0116 EN OUT0 VDD VSS / nand4
XI11 B net0105 VDD VSS / inverter
XI10 C net0116 VDD VSS / inverter
XI8 A net0158 VDD VSS / inverter
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG BL OUT SEL_B VDD VSS
*.PININFO BL:I SEL_B:I VDD:I VSS:I OUT:O
XI1 SEL_B net40 VDD VSS / inverter
MM1 BL net40 OUT VSS N_18 W=500.0n L=180.00n
MM0 BL SEL_B OUT VDD P_18 W=1.5u L=180.00n
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    YMUX
* View Name:    schematic
************************************************************************

.SUBCKT YMUX BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> Dout VDD VSS 
+ Ysel<0> Ysel<1> Ysel<2> Ysel<3> Ysel<4> Ysel<5> Ysel<6> Ysel<7>
*.PININFO BL<0>:I BL<1>:I BL<2>:I BL<3>:I BL<4>:I BL<5>:I BL<6>:I BL<7>:I 
*.PININFO Ysel<0>:I Ysel<1>:I Ysel<2>:I Ysel<3>:I Ysel<4>:I Ysel<5>:I 
*.PININFO Ysel<6>:I Ysel<7>:I Dout:O VDD:B VSS:B
XI15 BL<4> Dout Ysel<4> VDD VSS / TG
XI18 BL<7> Dout Ysel<7> VDD VSS / TG
XI19 BL<3> Dout Ysel<3> VDD VSS / TG
XI20 BL<2> Dout Ysel<2> VDD VSS / TG
XI21 BL<1> Dout Ysel<1> VDD VSS / TG
XI22 BL<0> Dout Ysel<0> VDD VSS / TG
XI16 BL<5> Dout Ysel<5> VDD VSS / TG
XI17 BL<6> Dout Ysel<6> VDD VSS / TG
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    precharge
* View Name:    schematic
************************************************************************

.SUBCKT precharge BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> 
+ BL<10> BL<11> BL<12> BL<13> BL<14> BL<15> VDD pre_b
*.PININFO BL<0>:I BL<1>:I BL<2>:I BL<3>:I BL<4>:I BL<5>:I BL<6>:I BL<7>:I 
*.PININFO BL<8>:I BL<9>:I BL<10>:I BL<11>:I BL<12>:I BL<13>:I BL<14>:I 
*.PININFO BL<15>:I VDD:I pre_b:I
MM8 BL<0> pre_b VDD VDD P_18 W=1.5u L=180n
MM9 BL<1> pre_b VDD VDD P_18 W=1.5u L=180n
MM10 BL<2> pre_b VDD VDD P_18 W=1.5u L=180n
MM11 BL<3> pre_b VDD VDD P_18 W=1.5u L=180n
MM12 BL<4> pre_b VDD VDD P_18 W=1.5u L=180n
MM13 BL<5> pre_b VDD VDD P_18 W=1.5u L=180n
MM14 BL<6> pre_b VDD VDD P_18 W=1.5u L=180n
MM15 BL<7> pre_b VDD VDD P_18 W=1.5u L=180n
MM7 BL<8> pre_b VDD VDD P_18 W=1.5u L=180n
MM6 BL<9> pre_b VDD VDD P_18 W=1.5u L=180n
MM5 BL<10> pre_b VDD VDD P_18 W=1.5u L=180n
MM4 BL<11> pre_b VDD VDD P_18 W=1.5u L=180n
MM3 BL<12> pre_b VDD VDD P_18 W=1.5u L=180n
MM2 BL<13> pre_b VDD VDD P_18 W=1.5u L=180n
MM1 BL<14> pre_b VDD VDD P_18 W=1.5u L=180n
MM0 BL<15> pre_b VDD VDD P_18 W=1.5u L=180n
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    ROM
* View Name:    schematic
************************************************************************

.SUBCKT ROM BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> 
+ BL<11> BL<12> BL<13> BL<14> BL<15> VSS WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> 
+ WL<6> WL<7> WL<8> WL<9> WL<10> WL<11> WL<12> WL<13> WL<14> WL<15> WL<16> 
+ WL<17> WL<18> WL<19> WL<20> WL<21> WL<22> WL<23> WL<24> WL<25> WL<26> WL<27> 
+ WL<28> WL<29> WL<30> WL<31> WL<32> WL<33> WL<34> WL<35> WL<36> WL<37> WL<38> 
+ WL<39> WL<40> WL<41> WL<42> WL<43> WL<44> WL<45> WL<46> WL<47> WL<48> WL<49> 
+ WL<50> WL<51> WL<52> WL<53> WL<54> WL<55> WL<56> WL<57> WL<58> WL<59> WL<60> 
+ WL<61> WL<62> WL<63>
*.PININFO VSS:I WL<0>:I WL<1>:I WL<2>:I WL<3>:I WL<4>:I WL<5>:I WL<6>:I 
*.PININFO WL<7>:I WL<8>:I WL<9>:I WL<10>:I WL<11>:I WL<12>:I WL<13>:I WL<14>:I 
*.PININFO WL<15>:I WL<16>:I WL<17>:I WL<18>:I WL<19>:I WL<20>:I WL<21>:I 
*.PININFO WL<22>:I WL<23>:I WL<24>:I WL<25>:I WL<26>:I WL<27>:I WL<28>:I 
*.PININFO WL<29>:I WL<30>:I WL<31>:I WL<32>:I WL<33>:I WL<34>:I WL<35>:I 
*.PININFO WL<36>:I WL<37>:I WL<38>:I WL<39>:I WL<40>:I WL<41>:I WL<42>:I 
*.PININFO WL<43>:I WL<44>:I WL<45>:I WL<46>:I WL<47>:I WL<48>:I WL<49>:I 
*.PININFO WL<50>:I WL<51>:I WL<52>:I WL<53>:I WL<54>:I WL<55>:I WL<56>:I 
*.PININFO WL<57>:I WL<58>:I WL<59>:I WL<60>:I WL<61>:I WL<62>:I WL<63>:I 
*.PININFO BL<0>:O BL<1>:O BL<2>:O BL<3>:O BL<4>:O BL<5>:O BL<6>:O BL<7>:O 
*.PININFO BL<8>:O BL<9>:O BL<10>:O BL<11>:O BL<12>:O BL<13>:O BL<14>:O BL<15>:O
MM1565 VSS WL<8> net1712 VSS N_18 W=470n L=180.00n
MM1564 VSS WL<8> BL<1> VSS N_18 W=470n L=180.00n
MM1562 VSS WL<9> net1720 VSS N_18 W=470n L=180.00n
MM1558 VSS WL<9> BL<12> VSS N_18 W=470n L=180.00n
MM1549 VSS WL<8> net1728 VSS N_18 W=470n L=180.00n
MM1546 VSS WL<11> net1732 VSS N_18 W=470n L=180.00n
MM1544 VSS WL<8> BL<3> VSS N_18 W=470n L=180.00n
MM1542 VSS WL<11> BL<10> VSS N_18 W=470n L=180.00n
MM1541 VSS WL<9> net1744 VSS N_18 W=470n L=180.00n
MM1540 VSS WL<11> net1748 VSS N_18 W=470n L=180.00n
MM1539 VSS WL<9> BL<0> VSS N_18 W=470n L=180.00n
MM1538 VSS WL<9> BL<2> VSS N_18 W=470n L=180.00n
MM1537 VSS WL<9> net1760 VSS N_18 W=470n L=180.00n
MM1536 VSS WL<9> net1764 VSS N_18 W=470n L=180.00n
MM1535 VSS WL<9> BL<4> VSS N_18 W=470n L=180.00n
MM1534 VSS WL<9> BL<6> VSS N_18 W=470n L=180.00n
MM1533 VSS WL<9> net1776 VSS N_18 W=470n L=180.00n
MM1532 VSS WL<9> net1780 VSS N_18 W=470n L=180.00n
MM1531 VSS WL<9> BL<8> VSS N_18 W=470n L=180.00n
MM1530 VSS WL<9> BL<10> VSS N_18 W=470n L=180.00n
MM1529 VSS WL<8> BL<5> VSS N_18 W=470n L=180.00n
MM1528 VSS WL<8> net1796 VSS N_18 W=470n L=180.00n
MM1527 VSS WL<8> net1800 VSS N_18 W=470n L=180.00n
MM1526 VSS WL<8> BL<7> VSS N_18 W=470n L=180.00n
MM1524 VSS WL<8> BL<9> VSS N_18 W=470n L=180.00n
MM1523 VSS WL<8> net1812 VSS N_18 W=470n L=180.00n
MM1522 VSS WL<12> net1816 VSS N_18 W=470n L=180.00n
MM1521 VSS WL<12> BL<1> VSS N_18 W=470n L=180.00n
MM1520 VSS WL<12> net1824 VSS N_18 W=470n L=180.00n
MM1519 VSS WL<12> BL<3> VSS N_18 W=470n L=180.00n
MM1518 VSS WL<12> BL<5> VSS N_18 W=470n L=180.00n
MM1517 VSS WL<12> net1836 VSS N_18 W=470n L=180.00n
MM1516 VSS WL<12> net1840 VSS N_18 W=470n L=180.00n
MM1515 VSS WL<12> BL<7> VSS N_18 W=470n L=180.00n
MM1514 VSS WL<12> BL<9> VSS N_18 W=470n L=180.00n
MM1513 VSS WL<12> net1852 VSS N_18 W=470n L=180.00n
MM1512 VSS WL<12> net1856 VSS N_18 W=470n L=180.00n
MM1511 VSS WL<12> BL<11> VSS N_18 W=470n L=180.00n
MM1510 VSS WL<12> BL<13> VSS N_18 W=470n L=180.00n
MM1509 VSS WL<12> net1868 VSS N_18 W=470n L=180.00n
MM1508 VSS WL<12> net1872 VSS N_18 W=470n L=180.00n
MM1507 VSS WL<12> BL<15> VSS N_18 W=470n L=180.00n
MM1103 VSS WL<1> BL<14> VSS N_18 W=470n L=180.00n
MM1127 VSS WL<3> BL<8> VSS N_18 W=470n L=180.00n
MM1128 VSS WL<3> net1888 VSS N_18 W=470n L=180.00n
MM1129 VSS WL<3> net1892 VSS N_18 W=470n L=180.00n
MM1130 VSS WL<3> BL<6> VSS N_18 W=470n L=180.00n
MM1131 VSS WL<3> BL<4> VSS N_18 W=470n L=180.00n
MM1132 VSS WL<3> net1904 VSS N_18 W=470n L=180.00n
MM1133 VSS WL<3> net1908 VSS N_18 W=470n L=180.00n
MM1134 VSS WL<3> BL<2> VSS N_18 W=470n L=180.00n
MM1135 VSS WL<3> BL<0> VSS N_18 W=470n L=180.00n
MM1136 VSS WL<3> net1920 VSS N_18 W=470n L=180.00n
MM1144 VSS WL<3> BL<12> VSS N_18 W=470n L=180.00n
MM1148 VSS WL<3> net1928 VSS N_18 W=470n L=180.00n
MM1166 VSS WL<2> BL<15> VSS N_18 W=470n L=180.00n
MM1167 VSS WL<2> net1936 VSS N_18 W=470n L=180.00n
MM1168 VSS WL<2> net1940 VSS N_18 W=470n L=180.00n
MM1169 VSS WL<2> BL<13> VSS N_18 W=470n L=180.00n
MM1170 VSS WL<2> BL<11> VSS N_18 W=470n L=180.00n
MM1171 VSS WL<2> net1952 VSS N_18 W=470n L=180.00n
MM1172 VSS WL<2> net1956 VSS N_18 W=470n L=180.00n
MM1173 VSS WL<2> BL<9> VSS N_18 W=470n L=180.00n
MM1174 VSS WL<2> BL<7> VSS N_18 W=470n L=180.00n
MM1175 VSS WL<2> net1968 VSS N_18 W=470n L=180.00n
MM1176 VSS WL<2> net1972 VSS N_18 W=470n L=180.00n
MM1177 VSS WL<2> BL<5> VSS N_18 W=470n L=180.00n
MM1178 VSS WL<2> BL<3> VSS N_18 W=470n L=180.00n
MM1179 VSS WL<2> net1984 VSS N_18 W=470n L=180.00n
MM1180 VSS WL<2> BL<1> VSS N_18 W=470n L=180.00n
MM1181 VSS WL<2> net1992 VSS N_18 W=470n L=180.00n
MM1106 VSS WL<1> net1996 VSS N_18 W=470n L=180.00n
MM1798 VSS WL<27> net2000 VSS N_18 W=470n L=180.00n
MM1780 VSS WL<26> BL<15> VSS N_18 W=470n L=180.00n
MM1779 VSS WL<26> net2008 VSS N_18 W=470n L=180.00n
MM1778 VSS WL<26> net2012 VSS N_18 W=470n L=180.00n
MM1777 VSS WL<26> BL<13> VSS N_18 W=470n L=180.00n
MM1776 VSS WL<26> BL<11> VSS N_18 W=470n L=180.00n
MM1775 VSS WL<26> net2024 VSS N_18 W=470n L=180.00n
MM1774 VSS WL<26> net2028 VSS N_18 W=470n L=180.00n
MM1773 VSS WL<26> BL<9> VSS N_18 W=470n L=180.00n
MM1772 VSS WL<26> BL<7> VSS N_18 W=470n L=180.00n
MM1771 VSS WL<26> net2040 VSS N_18 W=470n L=180.00n
MM1770 VSS WL<26> net2044 VSS N_18 W=470n L=180.00n
MM1769 VSS WL<26> BL<5> VSS N_18 W=470n L=180.00n
MM1768 VSS WL<26> BL<3> VSS N_18 W=470n L=180.00n
MM1767 VSS WL<26> net2056 VSS N_18 W=470n L=180.00n
MM1766 VSS WL<26> BL<1> VSS N_18 W=470n L=180.00n
MM1765 VSS WL<26> net2064 VSS N_18 W=470n L=180.00n
MM1753 VSS WL<25> net2068 VSS N_18 W=470n L=180.00n
MM1744 VSS WL<24> BL<15> VSS N_18 W=470n L=180.00n
MM1743 VSS WL<24> net2076 VSS N_18 W=470n L=180.00n
MM1742 VSS WL<30> net2080 VSS N_18 W=470n L=180.00n
MM1741 VSS WL<30> BL<1> VSS N_18 W=470n L=180.00n
MM1740 VSS WL<30> net2088 VSS N_18 W=470n L=180.00n
MM1739 VSS WL<30> BL<3> VSS N_18 W=470n L=180.00n
MM1738 VSS WL<30> BL<5> VSS N_18 W=470n L=180.00n
MM1737 VSS WL<30> net2100 VSS N_18 W=470n L=180.00n
MM1736 VSS WL<30> net2104 VSS N_18 W=470n L=180.00n
MM1735 VSS WL<30> BL<7> VSS N_18 W=470n L=180.00n
MM1734 VSS WL<30> BL<9> VSS N_18 W=470n L=180.00n
MM1733 VSS WL<30> net2116 VSS N_18 W=470n L=180.00n
MM1732 VSS WL<30> net2120 VSS N_18 W=470n L=180.00n
MM1731 VSS WL<30> BL<11> VSS N_18 W=470n L=180.00n
MM1730 VSS WL<30> BL<13> VSS N_18 W=470n L=180.00n
MM1729 VSS WL<30> net2132 VSS N_18 W=470n L=180.00n
MM1728 VSS WL<30> net2136 VSS N_18 W=470n L=180.00n
MM1727 VSS WL<30> BL<15> VSS N_18 W=470n L=180.00n
MM1719 VSS WL<25> net2144 VSS N_18 W=470n L=180.00n
MM1708 VSS WL<31> net2148 VSS N_18 W=470n L=180.00n
MM1704 VSS WL<31> BL<12> VSS N_18 W=470n L=180.00n
MM1696 VSS WL<31> net2156 VSS N_18 W=470n L=180.00n
MM1695 VSS WL<31> BL<0> VSS N_18 W=470n L=180.00n
MM1694 VSS WL<31> BL<2> VSS N_18 W=470n L=180.00n
MM1693 VSS WL<31> net2168 VSS N_18 W=470n L=180.00n
MM1692 VSS WL<31> net2172 VSS N_18 W=470n L=180.00n
MM1691 VSS WL<31> BL<4> VSS N_18 W=470n L=180.00n
MM1690 VSS WL<31> BL<6> VSS N_18 W=470n L=180.00n
MM1689 VSS WL<31> net2184 VSS N_18 W=470n L=180.00n
MM1688 VSS WL<31> net2188 VSS N_18 W=470n L=180.00n
MM1687 VSS WL<31> BL<8> VSS N_18 W=470n L=180.00n
MM1686 VSS WL<31> BL<10> VSS N_18 W=470n L=180.00n
MM1684 VSS WL<31> net2200 VSS N_18 W=470n L=180.00n
MM1683 VSS WL<31> net2204 VSS N_18 W=470n L=180.00n
MM1679 VSS WL<31> BL<14> VSS N_18 W=470n L=180.00n
MM1676 VSS WL<29> BL<14> VSS N_18 W=470n L=180.00n
MM1672 VSS WL<29> net2216 VSS N_18 W=470n L=180.00n
MM1671 VSS WL<29> net2220 VSS N_18 W=470n L=180.00n
MM1670 VSS WL<24> net2224 VSS N_18 W=470n L=180.00n
MM1668 VSS WL<29> BL<10> VSS N_18 W=470n L=180.00n
MM1667 VSS WL<29> BL<8> VSS N_18 W=470n L=180.00n
MM1666 VSS WL<29> net2236 VSS N_18 W=470n L=180.00n
MM1665 VSS WL<24> BL<13> VSS N_18 W=470n L=180.00n
MM1664 VSS WL<29> net2244 VSS N_18 W=470n L=180.00n
MM1663 VSS WL<24> BL<11> VSS N_18 W=470n L=180.00n
MM1662 VSS WL<29> BL<6> VSS N_18 W=470n L=180.00n
MM1661 VSS WL<29> BL<4> VSS N_18 W=470n L=180.00n
MM1660 VSS WL<29> net2260 VSS N_18 W=470n L=180.00n
MM1659 VSS WL<24> net2264 VSS N_18 W=470n L=180.00n
MM1658 VSS WL<29> net2268 VSS N_18 W=470n L=180.00n
MM1657 VSS WL<29> BL<2> VSS N_18 W=470n L=180.00n
MM1656 VSS WL<29> BL<0> VSS N_18 W=470n L=180.00n
MM1655 VSS WL<29> net2280 VSS N_18 W=470n L=180.00n
MM1647 VSS WL<27> BL<14> VSS N_18 W=470n L=180.00n
MM1646 VSS WL<29> BL<12> VSS N_18 W=470n L=180.00n
MM1642 VSS WL<29> net2292 VSS N_18 W=470n L=180.00n
MM1624 VSS WL<28> BL<15> VSS N_18 W=470n L=180.00n
MM1623 VSS WL<28> net2300 VSS N_18 W=470n L=180.00n
MM1622 VSS WL<28> net2304 VSS N_18 W=470n L=180.00n
MM1621 VSS WL<28> BL<13> VSS N_18 W=470n L=180.00n
MM1620 VSS WL<28> BL<11> VSS N_18 W=470n L=180.00n
MM1619 VSS WL<28> net2316 VSS N_18 W=470n L=180.00n
MM1618 VSS WL<28> net2320 VSS N_18 W=470n L=180.00n
MM1617 VSS WL<28> BL<9> VSS N_18 W=470n L=180.00n
MM1616 VSS WL<28> BL<7> VSS N_18 W=470n L=180.00n
MM1615 VSS WL<28> net2332 VSS N_18 W=470n L=180.00n
MM1614 VSS WL<28> net2336 VSS N_18 W=470n L=180.00n
MM1613 VSS WL<28> BL<5> VSS N_18 W=470n L=180.00n
MM1612 VSS WL<28> BL<3> VSS N_18 W=470n L=180.00n
MM1611 VSS WL<28> net2348 VSS N_18 W=470n L=180.00n
MM1610 VSS WL<28> BL<1> VSS N_18 W=470n L=180.00n
MM1609 VSS WL<28> net2356 VSS N_18 W=470n L=180.00n
MM1608 VSS WL<24> net2360 VSS N_18 W=470n L=180.00n
MM1607 VSS WL<24> BL<9> VSS N_18 W=470n L=180.00n
MM1605 VSS WL<24> BL<7> VSS N_18 W=470n L=180.00n
MM1604 VSS WL<24> net2372 VSS N_18 W=470n L=180.00n
MM1603 VSS WL<24> net2376 VSS N_18 W=470n L=180.00n
MM1602 VSS WL<24> BL<5> VSS N_18 W=470n L=180.00n
MM1601 VSS WL<25> BL<10> VSS N_18 W=470n L=180.00n
MM1600 VSS WL<25> BL<8> VSS N_18 W=470n L=180.00n
MM1599 VSS WL<25> net2392 VSS N_18 W=470n L=180.00n
MM1598 VSS WL<25> net2396 VSS N_18 W=470n L=180.00n
MM1597 VSS WL<25> BL<6> VSS N_18 W=470n L=180.00n
MM1596 VSS WL<25> BL<4> VSS N_18 W=470n L=180.00n
MM1595 VSS WL<25> net2408 VSS N_18 W=470n L=180.00n
MM1594 VSS WL<25> net2412 VSS N_18 W=470n L=180.00n
MM1593 VSS WL<25> BL<2> VSS N_18 W=470n L=180.00n
MM1592 VSS WL<25> BL<0> VSS N_18 W=470n L=180.00n
MM1591 VSS WL<27> net2424 VSS N_18 W=470n L=180.00n
MM1590 VSS WL<25> net2428 VSS N_18 W=470n L=180.00n
MM1589 VSS WL<27> BL<10> VSS N_18 W=470n L=180.00n
MM1587 VSS WL<24> BL<3> VSS N_18 W=470n L=180.00n
MM1585 VSS WL<27> net2440 VSS N_18 W=470n L=180.00n
MM1582 VSS WL<24> net2444 VSS N_18 W=470n L=180.00n
MM1573 VSS WL<25> BL<12> VSS N_18 W=470n L=180.00n
MM1569 VSS WL<25> net2452 VSS N_18 W=470n L=180.00n
MM1567 VSS WL<24> BL<1> VSS N_18 W=470n L=180.00n
MM1566 VSS WL<24> net2460 VSS N_18 W=470n L=180.00n
MM2077 VSS WL<16> net2464 VSS N_18 W=470n L=180.00n
MM2076 VSS WL<16> BL<1> VSS N_18 W=470n L=180.00n
MM2074 VSS WL<17> net2472 VSS N_18 W=470n L=180.00n
MM2070 VSS WL<17> BL<12> VSS N_18 W=470n L=180.00n
MM2061 VSS WL<16> net2480 VSS N_18 W=470n L=180.00n
MM2058 VSS WL<19> net2484 VSS N_18 W=470n L=180.00n
MM2056 VSS WL<16> BL<3> VSS N_18 W=470n L=180.00n
MM2054 VSS WL<19> BL<10> VSS N_18 W=470n L=180.00n
MM2053 VSS WL<17> net2496 VSS N_18 W=470n L=180.00n
MM2052 VSS WL<19> net2500 VSS N_18 W=470n L=180.00n
MM2051 VSS WL<17> BL<0> VSS N_18 W=470n L=180.00n
MM2050 VSS WL<17> BL<2> VSS N_18 W=470n L=180.00n
MM2049 VSS WL<17> net2512 VSS N_18 W=470n L=180.00n
MM2048 VSS WL<17> net2516 VSS N_18 W=470n L=180.00n
MM2047 VSS WL<17> BL<4> VSS N_18 W=470n L=180.00n
MM2046 VSS WL<17> BL<6> VSS N_18 W=470n L=180.00n
MM2045 VSS WL<17> net2528 VSS N_18 W=470n L=180.00n
MM2044 VSS WL<17> net2532 VSS N_18 W=470n L=180.00n
MM2043 VSS WL<17> BL<8> VSS N_18 W=470n L=180.00n
MM2042 VSS WL<17> BL<10> VSS N_18 W=470n L=180.00n
MM2041 VSS WL<16> BL<5> VSS N_18 W=470n L=180.00n
MM2040 VSS WL<16> net2548 VSS N_18 W=470n L=180.00n
MM2039 VSS WL<16> net2552 VSS N_18 W=470n L=180.00n
MM2038 VSS WL<16> BL<7> VSS N_18 W=470n L=180.00n
MM2036 VSS WL<16> BL<9> VSS N_18 W=470n L=180.00n
MM2035 VSS WL<16> net2564 VSS N_18 W=470n L=180.00n
MM2034 VSS WL<20> net02592 VSS N_18 W=470n L=180.00n
MM2033 VSS WL<20> BL<1> VSS N_18 W=470n L=180.00n
MM2032 VSS WL<20> net02600 VSS N_18 W=470n L=180.00n
MM2031 VSS WL<20> BL<3> VSS N_18 W=470n L=180.00n
MM2030 VSS WL<20> BL<5> VSS N_18 W=470n L=180.00n
MM2029 VSS WL<20> net02612 VSS N_18 W=470n L=180.00n
MM2028 VSS WL<20> net02616 VSS N_18 W=470n L=180.00n
MM2027 VSS WL<20> BL<7> VSS N_18 W=470n L=180.00n
MM2026 VSS WL<20> BL<9> VSS N_18 W=470n L=180.00n
MM2025 VSS WL<20> net02628 VSS N_18 W=470n L=180.00n
MM2024 VSS WL<20> net02632 VSS N_18 W=470n L=180.00n
MM2023 VSS WL<20> BL<11> VSS N_18 W=470n L=180.00n
MM2022 VSS WL<20> BL<13> VSS N_18 W=470n L=180.00n
MM2021 VSS WL<20> net02644 VSS N_18 W=470n L=180.00n
MM2020 VSS WL<20> net02641 VSS N_18 W=470n L=180.00n
MM2019 VSS WL<20> BL<15> VSS N_18 W=470n L=180.00n
MM2001 VSS WL<21> net2632 VSS N_18 W=470n L=180.00n
MM1997 VSS WL<21> BL<12> VSS N_18 W=470n L=180.00n
MM1996 VSS WL<19> BL<14> VSS N_18 W=470n L=180.00n
MM1988 VSS WL<21> net2644 VSS N_18 W=470n L=180.00n
MM1987 VSS WL<21> BL<0> VSS N_18 W=470n L=180.00n
MM1986 VSS WL<21> BL<2> VSS N_18 W=470n L=180.00n
MM1985 VSS WL<21> net2656 VSS N_18 W=470n L=180.00n
MM1984 VSS WL<16> net2660 VSS N_18 W=470n L=180.00n
MM1983 VSS WL<21> net2664 VSS N_18 W=470n L=180.00n
MM1982 VSS WL<21> BL<4> VSS N_18 W=470n L=180.00n
MM1981 VSS WL<21> BL<6> VSS N_18 W=470n L=180.00n
MM1980 VSS WL<16> BL<11> VSS N_18 W=470n L=180.00n
MM1979 VSS WL<21> net2680 VSS N_18 W=470n L=180.00n
MM1978 VSS WL<16> BL<13> VSS N_18 W=470n L=180.00n
MM1977 VSS WL<21> net2688 VSS N_18 W=470n L=180.00n
MM1976 VSS WL<21> BL<8> VSS N_18 W=470n L=180.00n
MM1975 VSS WL<21> BL<10> VSS N_18 W=470n L=180.00n
MM1973 VSS WL<16> net2700 VSS N_18 W=470n L=180.00n
MM1972 VSS WL<21> net2704 VSS N_18 W=470n L=180.00n
MM1971 VSS WL<21> net2708 VSS N_18 W=470n L=180.00n
MM1967 VSS WL<21> BL<14> VSS N_18 W=470n L=180.00n
MM1964 VSS WL<23> BL<14> VSS N_18 W=470n L=180.00n
MM1960 VSS WL<23> net2720 VSS N_18 W=470n L=180.00n
MM1959 VSS WL<23> net2724 VSS N_18 W=470n L=180.00n
MM1957 VSS WL<23> BL<10> VSS N_18 W=470n L=180.00n
MM1956 VSS WL<23> BL<8> VSS N_18 W=470n L=180.00n
MM1955 VSS WL<23> net2736 VSS N_18 W=470n L=180.00n
MM1954 VSS WL<23> net2740 VSS N_18 W=470n L=180.00n
MM1953 VSS WL<23> BL<6> VSS N_18 W=470n L=180.00n
MM1952 VSS WL<23> BL<4> VSS N_18 W=470n L=180.00n
MM1951 VSS WL<23> net2752 VSS N_18 W=470n L=180.00n
MM1950 VSS WL<23> net2756 VSS N_18 W=470n L=180.00n
MM1949 VSS WL<23> BL<2> VSS N_18 W=470n L=180.00n
MM1948 VSS WL<23> BL<0> VSS N_18 W=470n L=180.00n
MM1947 VSS WL<23> net2768 VSS N_18 W=470n L=180.00n
MM1939 VSS WL<23> BL<12> VSS N_18 W=470n L=180.00n
MM1935 VSS WL<23> net2776 VSS N_18 W=470n L=180.00n
MM1924 VSS WL<17> net2780 VSS N_18 W=470n L=180.00n
MM1916 VSS WL<22> BL<15> VSS N_18 W=470n L=180.00n
MM1915 VSS WL<22> net2788 VSS N_18 W=470n L=180.00n
MM1914 VSS WL<22> net2792 VSS N_18 W=470n L=180.00n
MM1913 VSS WL<22> BL<13> VSS N_18 W=470n L=180.00n
MM1912 VSS WL<22> BL<11> VSS N_18 W=470n L=180.00n
MM1911 VSS WL<22> net2804 VSS N_18 W=470n L=180.00n
MM1910 VSS WL<22> net2808 VSS N_18 W=470n L=180.00n
MM1909 VSS WL<22> BL<9> VSS N_18 W=470n L=180.00n
MM1908 VSS WL<22> BL<7> VSS N_18 W=470n L=180.00n
MM1907 VSS WL<22> net2820 VSS N_18 W=470n L=180.00n
MM1906 VSS WL<22> net2824 VSS N_18 W=470n L=180.00n
MM1905 VSS WL<22> BL<5> VSS N_18 W=470n L=180.00n
MM1904 VSS WL<22> BL<3> VSS N_18 W=470n L=180.00n
MM1903 VSS WL<22> net2836 VSS N_18 W=470n L=180.00n
MM1902 VSS WL<22> BL<1> VSS N_18 W=470n L=180.00n
MM1901 VSS WL<22> net2844 VSS N_18 W=470n L=180.00n
MM1900 VSS WL<16> net2848 VSS N_18 W=470n L=180.00n
MM1899 VSS WL<16> BL<15> VSS N_18 W=470n L=180.00n
MM1890 VSS WL<17> net2856 VSS N_18 W=470n L=180.00n
MM1878 VSS WL<18> net2860 VSS N_18 W=470n L=180.00n
MM1877 VSS WL<18> BL<1> VSS N_18 W=470n L=180.00n
MM1876 VSS WL<18> net2868 VSS N_18 W=470n L=180.00n
MM1875 VSS WL<18> BL<3> VSS N_18 W=470n L=180.00n
MM1874 VSS WL<18> BL<5> VSS N_18 W=470n L=180.00n
MM1873 VSS WL<18> net2880 VSS N_18 W=470n L=180.00n
MM1872 VSS WL<18> net2884 VSS N_18 W=470n L=180.00n
MM1871 VSS WL<18> BL<7> VSS N_18 W=470n L=180.00n
MM1870 VSS WL<18> BL<9> VSS N_18 W=470n L=180.00n
MM1869 VSS WL<18> net2896 VSS N_18 W=470n L=180.00n
MM1868 VSS WL<18> net2900 VSS N_18 W=470n L=180.00n
MM1867 VSS WL<18> BL<11> VSS N_18 W=470n L=180.00n
MM1866 VSS WL<18> BL<13> VSS N_18 W=470n L=180.00n
MM1865 VSS WL<18> net2912 VSS N_18 W=470n L=180.00n
MM1864 VSS WL<18> net2916 VSS N_18 W=470n L=180.00n
MM1863 VSS WL<18> BL<15> VSS N_18 W=470n L=180.00n
MM1845 VSS WL<19> net2924 VSS N_18 W=470n L=180.00n
MM1841 VSS WL<19> BL<12> VSS N_18 W=470n L=180.00n
MM1833 VSS WL<19> net2932 VSS N_18 W=470n L=180.00n
MM1832 VSS WL<19> BL<0> VSS N_18 W=470n L=180.00n
MM1831 VSS WL<19> BL<2> VSS N_18 W=470n L=180.00n
MM1830 VSS WL<19> net2944 VSS N_18 W=470n L=180.00n
MM1829 VSS WL<19> net2948 VSS N_18 W=470n L=180.00n
MM1828 VSS WL<19> BL<4> VSS N_18 W=470n L=180.00n
MM1827 VSS WL<19> BL<6> VSS N_18 W=470n L=180.00n
MM1826 VSS WL<19> net2960 VSS N_18 W=470n L=180.00n
MM1825 VSS WL<19> net2964 VSS N_18 W=470n L=180.00n
MM1824 VSS WL<19> BL<8> VSS N_18 W=470n L=180.00n
MM1823 VSS WL<17> BL<14> VSS N_18 W=470n L=180.00n
MM1820 VSS WL<25> BL<14> VSS N_18 W=470n L=180.00n
MM1819 VSS WL<27> BL<8> VSS N_18 W=470n L=180.00n
MM1818 VSS WL<27> net2984 VSS N_18 W=470n L=180.00n
MM1817 VSS WL<27> net2988 VSS N_18 W=470n L=180.00n
MM1816 VSS WL<27> BL<6> VSS N_18 W=470n L=180.00n
MM1815 VSS WL<27> BL<4> VSS N_18 W=470n L=180.00n
MM1814 VSS WL<27> net3000 VSS N_18 W=470n L=180.00n
MM1813 VSS WL<27> net3004 VSS N_18 W=470n L=180.00n
MM1812 VSS WL<27> BL<2> VSS N_18 W=470n L=180.00n
MM1811 VSS WL<27> BL<0> VSS N_18 W=470n L=180.00n
MM1810 VSS WL<27> net3016 VSS N_18 W=470n L=180.00n
MM1802 VSS WL<27> BL<12> VSS N_18 W=470n L=180.00n
MM1069 VSS WL<0> BL<15> VSS N_18 W=470n L=180.00n
MM1068 VSS WL<0> net3028 VSS N_18 W=470n L=180.00n
MM1182 VSS WL<6> net3032 VSS N_18 W=470n L=180.00n
MM1183 VSS WL<6> BL<1> VSS N_18 W=470n L=180.00n
MM1184 VSS WL<6> net3040 VSS N_18 W=470n L=180.00n
MM1185 VSS WL<6> BL<3> VSS N_18 W=470n L=180.00n
MM1186 VSS WL<6> BL<5> VSS N_18 W=470n L=180.00n
MM1187 VSS WL<6> net3052 VSS N_18 W=470n L=180.00n
MM1188 VSS WL<6> net3056 VSS N_18 W=470n L=180.00n
MM1189 VSS WL<6> BL<7> VSS N_18 W=470n L=180.00n
MM1190 VSS WL<6> BL<9> VSS N_18 W=470n L=180.00n
MM1191 VSS WL<6> net3068 VSS N_18 W=470n L=180.00n
MM1192 VSS WL<6> net3072 VSS N_18 W=470n L=180.00n
MM1193 VSS WL<6> BL<11> VSS N_18 W=470n L=180.00n
MM1194 VSS WL<6> BL<13> VSS N_18 W=470n L=180.00n
MM1195 VSS WL<6> net3084 VSS N_18 W=470n L=180.00n
MM1196 VSS WL<6> net3088 VSS N_18 W=470n L=180.00n
MM1197 VSS WL<6> BL<15> VSS N_18 W=470n L=180.00n
MM1105 VSS WL<1> net3096 VSS N_18 W=470n L=180.00n
MM1215 VSS WL<7> net3100 VSS N_18 W=470n L=180.00n
MM1219 VSS WL<7> BL<12> VSS N_18 W=470n L=180.00n
MM1227 VSS WL<7> net3108 VSS N_18 W=470n L=180.00n
MM1228 VSS WL<7> BL<0> VSS N_18 W=470n L=180.00n
MM1229 VSS WL<7> BL<2> VSS N_18 W=470n L=180.00n
MM1230 VSS WL<7> net3120 VSS N_18 W=470n L=180.00n
MM1231 VSS WL<7> net3124 VSS N_18 W=470n L=180.00n
MM1232 VSS WL<7> BL<4> VSS N_18 W=470n L=180.00n
MM1233 VSS WL<7> BL<6> VSS N_18 W=470n L=180.00n
MM1234 VSS WL<7> net3136 VSS N_18 W=470n L=180.00n
MM1235 VSS WL<7> net3140 VSS N_18 W=470n L=180.00n
MM1236 VSS WL<7> BL<8> VSS N_18 W=470n L=180.00n
MM1237 VSS WL<7> BL<10> VSS N_18 W=470n L=180.00n
MM1239 VSS WL<7> net3152 VSS N_18 W=470n L=180.00n
MM1240 VSS WL<7> net3156 VSS N_18 W=470n L=180.00n
MM1244 VSS WL<7> BL<14> VSS N_18 W=470n L=180.00n
MM1247 VSS WL<5> BL<14> VSS N_18 W=470n L=180.00n
MM1251 VSS WL<5> net3168 VSS N_18 W=470n L=180.00n
MM1252 VSS WL<5> net3172 VSS N_18 W=470n L=180.00n
MM1067 VSS WL<0> net3176 VSS N_18 W=470n L=180.00n
MM1254 VSS WL<5> BL<10> VSS N_18 W=470n L=180.00n
MM1255 VSS WL<5> BL<8> VSS N_18 W=470n L=180.00n
MM1256 VSS WL<5> net3188 VSS N_18 W=470n L=180.00n
MM1066 VSS WL<0> BL<13> VSS N_18 W=470n L=180.00n
MM1257 VSS WL<5> net3196 VSS N_18 W=470n L=180.00n
MM1065 VSS WL<0> BL<11> VSS N_18 W=470n L=180.00n
MM1258 VSS WL<5> BL<6> VSS N_18 W=470n L=180.00n
MM1259 VSS WL<5> BL<4> VSS N_18 W=470n L=180.00n
MM1260 VSS WL<5> net3212 VSS N_18 W=470n L=180.00n
MM1064 VSS WL<0> net3216 VSS N_18 W=470n L=180.00n
MM1261 VSS WL<5> net3220 VSS N_18 W=470n L=180.00n
MM1262 VSS WL<5> BL<2> VSS N_18 W=470n L=180.00n
MM1263 VSS WL<5> BL<0> VSS N_18 W=470n L=180.00n
MM1264 VSS WL<5> net3232 VSS N_18 W=470n L=180.00n
MM1119 VSS WL<3> BL<14> VSS N_18 W=470n L=180.00n
MM1272 VSS WL<5> BL<12> VSS N_18 W=470n L=180.00n
MM1276 VSS WL<5> net3244 VSS N_18 W=470n L=180.00n
MM1294 VSS WL<4> BL<15> VSS N_18 W=470n L=180.00n
MM1295 VSS WL<4> net3252 VSS N_18 W=470n L=180.00n
MM1296 VSS WL<4> net3256 VSS N_18 W=470n L=180.00n
MM1297 VSS WL<4> BL<13> VSS N_18 W=470n L=180.00n
MM1298 VSS WL<4> BL<11> VSS N_18 W=470n L=180.00n
MM1299 VSS WL<4> net3268 VSS N_18 W=470n L=180.00n
MM1300 VSS WL<4> net3272 VSS N_18 W=470n L=180.00n
MM1301 VSS WL<4> BL<9> VSS N_18 W=470n L=180.00n
MM1302 VSS WL<4> BL<7> VSS N_18 W=470n L=180.00n
MM1303 VSS WL<4> net3284 VSS N_18 W=470n L=180.00n
MM1304 VSS WL<4> net3288 VSS N_18 W=470n L=180.00n
MM1305 VSS WL<4> BL<5> VSS N_18 W=470n L=180.00n
MM1306 VSS WL<4> BL<3> VSS N_18 W=470n L=180.00n
MM1307 VSS WL<4> net3300 VSS N_18 W=470n L=180.00n
MM1308 VSS WL<4> BL<1> VSS N_18 W=470n L=180.00n
MM1309 VSS WL<4> net3308 VSS N_18 W=470n L=180.00n
MM1311 VSS WL<9> BL<14> VSS N_18 W=470n L=180.00n
MM1312 VSS WL<11> BL<8> VSS N_18 W=470n L=180.00n
MM1313 VSS WL<11> net3320 VSS N_18 W=470n L=180.00n
MM1314 VSS WL<11> net3324 VSS N_18 W=470n L=180.00n
MM1315 VSS WL<11> BL<6> VSS N_18 W=470n L=180.00n
MM1316 VSS WL<11> BL<4> VSS N_18 W=470n L=180.00n
MM1063 VSS WL<0> net3336 VSS N_18 W=470n L=180.00n
MM1062 VSS WL<0> BL<9> VSS N_18 W=470n L=180.00n
MM1061 VSS WL<0> BL<7> VSS N_18 W=470n L=180.00n
MM1060 VSS WL<0> net3348 VSS N_18 W=470n L=180.00n
MM1317 VSS WL<11> net3352 VSS N_18 W=470n L=180.00n
MM1318 VSS WL<11> net3356 VSS N_18 W=470n L=180.00n
MM1059 VSS WL<0> net3360 VSS N_18 W=470n L=180.00n
MM1058 VSS WL<0> BL<5> VSS N_18 W=470n L=180.00n
MM1319 VSS WL<11> BL<2> VSS N_18 W=470n L=180.00n
MM1320 VSS WL<11> BL<0> VSS N_18 W=470n L=180.00n
MM1107 VSS WL<1> BL<10> VSS N_18 W=470n L=180.00n
MM1108 VSS WL<1> BL<8> VSS N_18 W=470n L=180.00n
MM1109 VSS WL<1> net3384 VSS N_18 W=470n L=180.00n
MM1110 VSS WL<1> net3388 VSS N_18 W=470n L=180.00n
MM1111 VSS WL<1> BL<6> VSS N_18 W=470n L=180.00n
MM1112 VSS WL<1> BL<4> VSS N_18 W=470n L=180.00n
MM1113 VSS WL<1> net3400 VSS N_18 W=470n L=180.00n
MM1114 VSS WL<1> net3404 VSS N_18 W=470n L=180.00n
MM1115 VSS WL<1> BL<2> VSS N_18 W=470n L=180.00n
MM1116 VSS WL<1> BL<0> VSS N_18 W=470n L=180.00n
MM1123 VSS WL<3> net3416 VSS N_18 W=470n L=180.00n
MM1117 VSS WL<1> net3420 VSS N_18 W=470n L=180.00n
MM1126 VSS WL<3> BL<10> VSS N_18 W=470n L=180.00n
MM1057 VSS WL<0> BL<3> VSS N_18 W=470n L=180.00n
MM1321 VSS WL<11> net3432 VSS N_18 W=470n L=180.00n
MM1124 VSS WL<3> net3436 VSS N_18 W=470n L=180.00n
MM2136 VSS WL<52> BL<15> VSS N_18 W=470n L=180.00n
MM2135 VSS WL<52> net3444 VSS N_18 W=470n L=180.00n
MM2134 VSS WL<52> net3448 VSS N_18 W=470n L=180.00n
MM2133 VSS WL<52> BL<13> VSS N_18 W=470n L=180.00n
MM2132 VSS WL<52> BL<11> VSS N_18 W=470n L=180.00n
MM2131 VSS WL<52> net3460 VSS N_18 W=470n L=180.00n
MM2130 VSS WL<52> net3464 VSS N_18 W=470n L=180.00n
MM2129 VSS WL<52> BL<9> VSS N_18 W=470n L=180.00n
MM2128 VSS WL<52> BL<7> VSS N_18 W=470n L=180.00n
MM2127 VSS WL<52> net3476 VSS N_18 W=470n L=180.00n
MM2126 VSS WL<52> net3480 VSS N_18 W=470n L=180.00n
MM2125 VSS WL<52> BL<5> VSS N_18 W=470n L=180.00n
MM2124 VSS WL<52> BL<3> VSS N_18 W=470n L=180.00n
MM2123 VSS WL<52> net3492 VSS N_18 W=470n L=180.00n
MM2122 VSS WL<52> BL<1> VSS N_18 W=470n L=180.00n
MM2121 VSS WL<52> net3500 VSS N_18 W=470n L=180.00n
MM2120 VSS WL<48> net3504 VSS N_18 W=470n L=180.00n
MM2119 VSS WL<48> BL<9> VSS N_18 W=470n L=180.00n
MM2117 VSS WL<48> BL<7> VSS N_18 W=470n L=180.00n
MM2116 VSS WL<48> net3516 VSS N_18 W=470n L=180.00n
MM2115 VSS WL<48> net3520 VSS N_18 W=470n L=180.00n
MM2114 VSS WL<48> BL<5> VSS N_18 W=470n L=180.00n
MM2113 VSS WL<49> BL<10> VSS N_18 W=470n L=180.00n
MM2112 VSS WL<49> BL<8> VSS N_18 W=470n L=180.00n
MM2111 VSS WL<49> net3536 VSS N_18 W=470n L=180.00n
MM2110 VSS WL<49> net3540 VSS N_18 W=470n L=180.00n
MM2109 VSS WL<49> BL<6> VSS N_18 W=470n L=180.00n
MM2108 VSS WL<49> BL<4> VSS N_18 W=470n L=180.00n
MM2107 VSS WL<49> net3552 VSS N_18 W=470n L=180.00n
MM2106 VSS WL<49> net3556 VSS N_18 W=470n L=180.00n
MM2105 VSS WL<49> BL<2> VSS N_18 W=470n L=180.00n
MM2104 VSS WL<49> BL<0> VSS N_18 W=470n L=180.00n
MM2103 VSS WL<51> net3568 VSS N_18 W=470n L=180.00n
MM2102 VSS WL<49> net3572 VSS N_18 W=470n L=180.00n
MM2101 VSS WL<51> BL<10> VSS N_18 W=470n L=180.00n
MM2099 VSS WL<48> BL<3> VSS N_18 W=470n L=180.00n
MM2097 VSS WL<51> net3584 VSS N_18 W=470n L=180.00n
MM2094 VSS WL<48> net3588 VSS N_18 W=470n L=180.00n
MM2085 VSS WL<49> BL<12> VSS N_18 W=470n L=180.00n
MM2081 VSS WL<49> net3596 VSS N_18 W=470n L=180.00n
MM2079 VSS WL<48> BL<1> VSS N_18 W=470n L=180.00n
MM2078 VSS WL<48> net3604 VSS N_18 W=470n L=180.00n
MM2495 VSS WL<61> net3608 VSS N_18 W=470n L=180.00n
MM2494 VSS WL<61> BL<4> VSS N_18 W=470n L=180.00n
MM2493 VSS WL<61> BL<6> VSS N_18 W=470n L=180.00n
MM2492 VSS WL<56> BL<11> VSS N_18 W=470n L=180.00n
MM2491 VSS WL<61> net3624 VSS N_18 W=470n L=180.00n
MM2490 VSS WL<56> BL<13> VSS N_18 W=470n L=180.00n
MM2489 VSS WL<61> net3632 VSS N_18 W=470n L=180.00n
MM2488 VSS WL<61> BL<8> VSS N_18 W=470n L=180.00n
MM2487 VSS WL<61> BL<10> VSS N_18 W=470n L=180.00n
MM2485 VSS WL<56> net3644 VSS N_18 W=470n L=180.00n
MM2484 VSS WL<61> net3648 VSS N_18 W=470n L=180.00n
MM2483 VSS WL<61> net3652 VSS N_18 W=470n L=180.00n
MM2479 VSS WL<61> BL<14> VSS N_18 W=470n L=180.00n
MM2476 VSS WL<63> BL<14> VSS N_18 W=470n L=180.00n
MM2472 VSS WL<63> net3664 VSS N_18 W=470n L=180.00n
MM2471 VSS WL<63> net3668 VSS N_18 W=470n L=180.00n
MM2469 VSS WL<63> BL<10> VSS N_18 W=470n L=180.00n
MM2468 VSS WL<63> BL<8> VSS N_18 W=470n L=180.00n
MM2467 VSS WL<63> net3680 VSS N_18 W=470n L=180.00n
MM2466 VSS WL<63> net3684 VSS N_18 W=470n L=180.00n
MM2465 VSS WL<63> BL<6> VSS N_18 W=470n L=180.00n
MM2464 VSS WL<63> BL<4> VSS N_18 W=470n L=180.00n
MM2463 VSS WL<63> net3696 VSS N_18 W=470n L=180.00n
MM2462 VSS WL<63> net3700 VSS N_18 W=470n L=180.00n
MM2461 VSS WL<63> BL<2> VSS N_18 W=470n L=180.00n
MM2460 VSS WL<63> BL<0> VSS N_18 W=470n L=180.00n
MM2459 VSS WL<63> net3712 VSS N_18 W=470n L=180.00n
MM2451 VSS WL<63> BL<12> VSS N_18 W=470n L=180.00n
MM2447 VSS WL<63> net3720 VSS N_18 W=470n L=180.00n
MM2436 VSS WL<57> net3724 VSS N_18 W=470n L=180.00n
MM2428 VSS WL<62> BL<15> VSS N_18 W=470n L=180.00n
MM2427 VSS WL<62> net3732 VSS N_18 W=470n L=180.00n
MM2426 VSS WL<62> net3736 VSS N_18 W=470n L=180.00n
MM2425 VSS WL<62> BL<13> VSS N_18 W=470n L=180.00n
MM2424 VSS WL<62> BL<11> VSS N_18 W=470n L=180.00n
MM2423 VSS WL<62> net3748 VSS N_18 W=470n L=180.00n
MM2422 VSS WL<62> net3752 VSS N_18 W=470n L=180.00n
MM2421 VSS WL<62> BL<9> VSS N_18 W=470n L=180.00n
MM2420 VSS WL<62> BL<7> VSS N_18 W=470n L=180.00n
MM2419 VSS WL<62> net3764 VSS N_18 W=470n L=180.00n
MM2418 VSS WL<62> net3768 VSS N_18 W=470n L=180.00n
MM2417 VSS WL<62> BL<5> VSS N_18 W=470n L=180.00n
MM2416 VSS WL<62> BL<3> VSS N_18 W=470n L=180.00n
MM2415 VSS WL<62> net3780 VSS N_18 W=470n L=180.00n
MM2414 VSS WL<62> BL<1> VSS N_18 W=470n L=180.00n
MM2413 VSS WL<62> net3788 VSS N_18 W=470n L=180.00n
MM2412 VSS WL<56> net3792 VSS N_18 W=470n L=180.00n
MM2411 VSS WL<56> BL<15> VSS N_18 W=470n L=180.00n
MM2402 VSS WL<57> net3800 VSS N_18 W=470n L=180.00n
MM2390 VSS WL<58> net3804 VSS N_18 W=470n L=180.00n
MM2389 VSS WL<58> BL<1> VSS N_18 W=470n L=180.00n
MM2388 VSS WL<58> net3812 VSS N_18 W=470n L=180.00n
MM2387 VSS WL<58> BL<3> VSS N_18 W=470n L=180.00n
MM2386 VSS WL<58> BL<5> VSS N_18 W=470n L=180.00n
MM2385 VSS WL<58> net3824 VSS N_18 W=470n L=180.00n
MM2384 VSS WL<58> net3828 VSS N_18 W=470n L=180.00n
MM2383 VSS WL<58> BL<7> VSS N_18 W=470n L=180.00n
MM2382 VSS WL<58> BL<9> VSS N_18 W=470n L=180.00n
MM2381 VSS WL<58> net3840 VSS N_18 W=470n L=180.00n
MM2380 VSS WL<58> net3844 VSS N_18 W=470n L=180.00n
MM2379 VSS WL<58> BL<11> VSS N_18 W=470n L=180.00n
MM2378 VSS WL<58> BL<13> VSS N_18 W=470n L=180.00n
MM2377 VSS WL<58> net3856 VSS N_18 W=470n L=180.00n
MM2376 VSS WL<58> net3860 VSS N_18 W=470n L=180.00n
MM2375 VSS WL<58> BL<15> VSS N_18 W=470n L=180.00n
MM2357 VSS WL<59> net3868 VSS N_18 W=470n L=180.00n
MM2353 VSS WL<59> BL<12> VSS N_18 W=470n L=180.00n
MM2345 VSS WL<59> net3876 VSS N_18 W=470n L=180.00n
MM2344 VSS WL<59> BL<0> VSS N_18 W=470n L=180.00n
MM2343 VSS WL<59> BL<2> VSS N_18 W=470n L=180.00n
MM2342 VSS WL<59> net3888 VSS N_18 W=470n L=180.00n
MM2341 VSS WL<59> net3892 VSS N_18 W=470n L=180.00n
MM2340 VSS WL<59> BL<4> VSS N_18 W=470n L=180.00n
MM2339 VSS WL<59> BL<6> VSS N_18 W=470n L=180.00n
MM2338 VSS WL<59> net3904 VSS N_18 W=470n L=180.00n
MM2337 VSS WL<59> net3908 VSS N_18 W=470n L=180.00n
MM2336 VSS WL<59> BL<8> VSS N_18 W=470n L=180.00n
MM2335 VSS WL<57> BL<14> VSS N_18 W=470n L=180.00n
MM2332 VSS WL<49> BL<14> VSS N_18 W=470n L=180.00n
MM2331 VSS WL<51> BL<8> VSS N_18 W=470n L=180.00n
MM2330 VSS WL<51> net3928 VSS N_18 W=470n L=180.00n
MM2329 VSS WL<51> net3932 VSS N_18 W=470n L=180.00n
MM2328 VSS WL<51> BL<6> VSS N_18 W=470n L=180.00n
MM2327 VSS WL<51> BL<4> VSS N_18 W=470n L=180.00n
MM2326 VSS WL<51> net3944 VSS N_18 W=470n L=180.00n
MM2325 VSS WL<51> net3948 VSS N_18 W=470n L=180.00n
MM2324 VSS WL<51> BL<2> VSS N_18 W=470n L=180.00n
MM2323 VSS WL<51> BL<0> VSS N_18 W=470n L=180.00n
MM2322 VSS WL<51> net3960 VSS N_18 W=470n L=180.00n
MM2314 VSS WL<51> BL<12> VSS N_18 W=470n L=180.00n
MM2310 VSS WL<51> net3968 VSS N_18 W=470n L=180.00n
MM2292 VSS WL<50> BL<15> VSS N_18 W=470n L=180.00n
MM2291 VSS WL<50> net3976 VSS N_18 W=470n L=180.00n
MM2290 VSS WL<50> net3980 VSS N_18 W=470n L=180.00n
MM2289 VSS WL<50> BL<13> VSS N_18 W=470n L=180.00n
MM2288 VSS WL<50> BL<11> VSS N_18 W=470n L=180.00n
MM2287 VSS WL<50> net3992 VSS N_18 W=470n L=180.00n
MM2286 VSS WL<50> net3996 VSS N_18 W=470n L=180.00n
MM2285 VSS WL<50> BL<9> VSS N_18 W=470n L=180.00n
MM2284 VSS WL<50> BL<7> VSS N_18 W=470n L=180.00n
MM2283 VSS WL<50> net4008 VSS N_18 W=470n L=180.00n
MM2282 VSS WL<50> net4012 VSS N_18 W=470n L=180.00n
MM2281 VSS WL<50> BL<5> VSS N_18 W=470n L=180.00n
MM2280 VSS WL<50> BL<3> VSS N_18 W=470n L=180.00n
MM2279 VSS WL<50> net4024 VSS N_18 W=470n L=180.00n
MM2278 VSS WL<50> BL<1> VSS N_18 W=470n L=180.00n
MM2277 VSS WL<50> net4032 VSS N_18 W=470n L=180.00n
MM2265 VSS WL<49> net4036 VSS N_18 W=470n L=180.00n
MM2256 VSS WL<48> BL<15> VSS N_18 W=470n L=180.00n
MM2255 VSS WL<48> net4044 VSS N_18 W=470n L=180.00n
MM2254 VSS WL<54> net4048 VSS N_18 W=470n L=180.00n
MM2253 VSS WL<54> BL<1> VSS N_18 W=470n L=180.00n
MM2252 VSS WL<54> net4056 VSS N_18 W=470n L=180.00n
MM2251 VSS WL<54> BL<3> VSS N_18 W=470n L=180.00n
MM2250 VSS WL<54> BL<5> VSS N_18 W=470n L=180.00n
MM2249 VSS WL<54> net4068 VSS N_18 W=470n L=180.00n
MM2248 VSS WL<54> net4072 VSS N_18 W=470n L=180.00n
MM2247 VSS WL<54> BL<7> VSS N_18 W=470n L=180.00n
MM2246 VSS WL<54> BL<9> VSS N_18 W=470n L=180.00n
MM2245 VSS WL<54> net4084 VSS N_18 W=470n L=180.00n
MM2244 VSS WL<54> net4088 VSS N_18 W=470n L=180.00n
MM2243 VSS WL<54> BL<11> VSS N_18 W=470n L=180.00n
MM2242 VSS WL<54> BL<13> VSS N_18 W=470n L=180.00n
MM2241 VSS WL<54> net4100 VSS N_18 W=470n L=180.00n
MM2240 VSS WL<54> net4104 VSS N_18 W=470n L=180.00n
MM2239 VSS WL<54> BL<15> VSS N_18 W=470n L=180.00n
MM2231 VSS WL<49> net4112 VSS N_18 W=470n L=180.00n
MM2220 VSS WL<55> net4116 VSS N_18 W=470n L=180.00n
MM2216 VSS WL<55> BL<12> VSS N_18 W=470n L=180.00n
MM2208 VSS WL<55> net4124 VSS N_18 W=470n L=180.00n
MM2207 VSS WL<55> BL<0> VSS N_18 W=470n L=180.00n
MM2206 VSS WL<55> BL<2> VSS N_18 W=470n L=180.00n
MM2205 VSS WL<55> net4136 VSS N_18 W=470n L=180.00n
MM2204 VSS WL<55> net4140 VSS N_18 W=470n L=180.00n
MM2203 VSS WL<55> BL<4> VSS N_18 W=470n L=180.00n
MM2202 VSS WL<55> BL<6> VSS N_18 W=470n L=180.00n
MM2201 VSS WL<55> net4152 VSS N_18 W=470n L=180.00n
MM2200 VSS WL<55> net4156 VSS N_18 W=470n L=180.00n
MM2199 VSS WL<55> BL<8> VSS N_18 W=470n L=180.00n
MM2198 VSS WL<55> BL<10> VSS N_18 W=470n L=180.00n
MM2196 VSS WL<55> net4168 VSS N_18 W=470n L=180.00n
MM2195 VSS WL<55> net4172 VSS N_18 W=470n L=180.00n
MM2191 VSS WL<55> BL<14> VSS N_18 W=470n L=180.00n
MM2188 VSS WL<53> BL<14> VSS N_18 W=470n L=180.00n
MM2184 VSS WL<53> net4184 VSS N_18 W=470n L=180.00n
MM2183 VSS WL<53> net4188 VSS N_18 W=470n L=180.00n
MM2182 VSS WL<48> net4192 VSS N_18 W=470n L=180.00n
MM2180 VSS WL<53> BL<10> VSS N_18 W=470n L=180.00n
MM2179 VSS WL<53> BL<8> VSS N_18 W=470n L=180.00n
MM2178 VSS WL<53> net4204 VSS N_18 W=470n L=180.00n
MM2177 VSS WL<48> BL<13> VSS N_18 W=470n L=180.00n
MM2176 VSS WL<53> net4212 VSS N_18 W=470n L=180.00n
MM2175 VSS WL<48> BL<11> VSS N_18 W=470n L=180.00n
MM2174 VSS WL<53> BL<6> VSS N_18 W=470n L=180.00n
MM2173 VSS WL<53> BL<4> VSS N_18 W=470n L=180.00n
MM2172 VSS WL<53> net4228 VSS N_18 W=470n L=180.00n
MM2171 VSS WL<48> net4232 VSS N_18 W=470n L=180.00n
MM2170 VSS WL<53> net4236 VSS N_18 W=470n L=180.00n
MM2169 VSS WL<53> BL<2> VSS N_18 W=470n L=180.00n
MM2168 VSS WL<53> BL<0> VSS N_18 W=470n L=180.00n
MM2167 VSS WL<53> net4248 VSS N_18 W=470n L=180.00n
MM2159 VSS WL<51> BL<14> VSS N_18 W=470n L=180.00n
MM2158 VSS WL<53> BL<12> VSS N_18 W=470n L=180.00n
MM2154 VSS WL<53> net4260 VSS N_18 W=470n L=180.00n
MM1056 VSS WL<0> net4264 VSS N_18 W=470n L=180.00n
MM2914 VSS WL<33> net4268 VSS N_18 W=470n L=180.00n
MM2902 VSS WL<34> net4272 VSS N_18 W=470n L=180.00n
MM2901 VSS WL<34> BL<1> VSS N_18 W=470n L=180.00n
MM2900 VSS WL<34> net4280 VSS N_18 W=470n L=180.00n
MM2899 VSS WL<34> BL<3> VSS N_18 W=470n L=180.00n
MM2898 VSS WL<34> BL<5> VSS N_18 W=470n L=180.00n
MM2897 VSS WL<34> net4292 VSS N_18 W=470n L=180.00n
MM2896 VSS WL<34> net4296 VSS N_18 W=470n L=180.00n
MM2895 VSS WL<34> BL<7> VSS N_18 W=470n L=180.00n
MM2894 VSS WL<34> BL<9> VSS N_18 W=470n L=180.00n
MM2893 VSS WL<34> net4308 VSS N_18 W=470n L=180.00n
MM2892 VSS WL<34> net4312 VSS N_18 W=470n L=180.00n
MM2891 VSS WL<34> BL<11> VSS N_18 W=470n L=180.00n
MM2890 VSS WL<34> BL<13> VSS N_18 W=470n L=180.00n
MM2889 VSS WL<34> net4324 VSS N_18 W=470n L=180.00n
MM2888 VSS WL<34> net4328 VSS N_18 W=470n L=180.00n
MM2887 VSS WL<34> BL<15> VSS N_18 W=470n L=180.00n
MM2869 VSS WL<35> net4336 VSS N_18 W=470n L=180.00n
MM2865 VSS WL<35> BL<12> VSS N_18 W=470n L=180.00n
MM2857 VSS WL<35> net4344 VSS N_18 W=470n L=180.00n
MM2856 VSS WL<35> BL<0> VSS N_18 W=470n L=180.00n
MM2855 VSS WL<35> BL<2> VSS N_18 W=470n L=180.00n
MM2854 VSS WL<35> net4356 VSS N_18 W=470n L=180.00n
MM2853 VSS WL<35> net4360 VSS N_18 W=470n L=180.00n
MM2852 VSS WL<35> BL<4> VSS N_18 W=470n L=180.00n
MM2851 VSS WL<35> BL<6> VSS N_18 W=470n L=180.00n
MM2850 VSS WL<35> net4372 VSS N_18 W=470n L=180.00n
MM2849 VSS WL<35> net4376 VSS N_18 W=470n L=180.00n
MM2848 VSS WL<35> BL<8> VSS N_18 W=470n L=180.00n
MM2847 VSS WL<33> BL<14> VSS N_18 W=470n L=180.00n
MM2844 VSS WL<41> BL<14> VSS N_18 W=470n L=180.00n
MM2843 VSS WL<43> BL<8> VSS N_18 W=470n L=180.00n
MM2842 VSS WL<43> net4396 VSS N_18 W=470n L=180.00n
MM2841 VSS WL<43> net4400 VSS N_18 W=470n L=180.00n
MM2840 VSS WL<43> BL<6> VSS N_18 W=470n L=180.00n
MM2839 VSS WL<43> BL<4> VSS N_18 W=470n L=180.00n
MM2838 VSS WL<43> net4412 VSS N_18 W=470n L=180.00n
MM2837 VSS WL<43> net4416 VSS N_18 W=470n L=180.00n
MM2836 VSS WL<43> BL<2> VSS N_18 W=470n L=180.00n
MM2835 VSS WL<43> BL<0> VSS N_18 W=470n L=180.00n
MM2834 VSS WL<43> net4428 VSS N_18 W=470n L=180.00n
MM2826 VSS WL<43> BL<12> VSS N_18 W=470n L=180.00n
MM2822 VSS WL<43> net4436 VSS N_18 W=470n L=180.00n
MM2804 VSS WL<42> BL<15> VSS N_18 W=470n L=180.00n
MM2803 VSS WL<42> net4444 VSS N_18 W=470n L=180.00n
MM2802 VSS WL<42> net4448 VSS N_18 W=470n L=180.00n
MM2801 VSS WL<42> BL<13> VSS N_18 W=470n L=180.00n
MM2800 VSS WL<42> BL<11> VSS N_18 W=470n L=180.00n
MM2799 VSS WL<42> net4460 VSS N_18 W=470n L=180.00n
MM2798 VSS WL<42> net4464 VSS N_18 W=470n L=180.00n
MM2797 VSS WL<42> BL<9> VSS N_18 W=470n L=180.00n
MM2796 VSS WL<42> BL<7> VSS N_18 W=470n L=180.00n
MM2795 VSS WL<42> net4476 VSS N_18 W=470n L=180.00n
MM2794 VSS WL<42> net4480 VSS N_18 W=470n L=180.00n
MM2793 VSS WL<42> BL<5> VSS N_18 W=470n L=180.00n
MM2792 VSS WL<42> BL<3> VSS N_18 W=470n L=180.00n
MM2791 VSS WL<42> net4492 VSS N_18 W=470n L=180.00n
MM2790 VSS WL<42> BL<1> VSS N_18 W=470n L=180.00n
MM2789 VSS WL<42> net4500 VSS N_18 W=470n L=180.00n
MM2777 VSS WL<41> net4504 VSS N_18 W=470n L=180.00n
MM2768 VSS WL<40> BL<15> VSS N_18 W=470n L=180.00n
MM2767 VSS WL<40> net4512 VSS N_18 W=470n L=180.00n
MM2766 VSS WL<46> net4516 VSS N_18 W=470n L=180.00n
MM2765 VSS WL<46> BL<1> VSS N_18 W=470n L=180.00n
MM2764 VSS WL<46> net4524 VSS N_18 W=470n L=180.00n
MM2763 VSS WL<46> BL<3> VSS N_18 W=470n L=180.00n
MM2762 VSS WL<46> BL<5> VSS N_18 W=470n L=180.00n
MM2761 VSS WL<46> net4536 VSS N_18 W=470n L=180.00n
MM2760 VSS WL<46> net4540 VSS N_18 W=470n L=180.00n
MM2759 VSS WL<46> BL<7> VSS N_18 W=470n L=180.00n
MM2758 VSS WL<46> BL<9> VSS N_18 W=470n L=180.00n
MM2757 VSS WL<46> net4552 VSS N_18 W=470n L=180.00n
MM2756 VSS WL<46> net4556 VSS N_18 W=470n L=180.00n
MM2755 VSS WL<46> BL<11> VSS N_18 W=470n L=180.00n
MM2754 VSS WL<46> BL<13> VSS N_18 W=470n L=180.00n
MM2753 VSS WL<46> net4568 VSS N_18 W=470n L=180.00n
MM2752 VSS WL<46> net4572 VSS N_18 W=470n L=180.00n
MM2751 VSS WL<46> BL<15> VSS N_18 W=470n L=180.00n
MM2743 VSS WL<41> net4580 VSS N_18 W=470n L=180.00n
MM2732 VSS WL<47> net4584 VSS N_18 W=470n L=180.00n
MM2728 VSS WL<47> BL<12> VSS N_18 W=470n L=180.00n
MM2720 VSS WL<47> net4592 VSS N_18 W=470n L=180.00n
MM2719 VSS WL<47> BL<0> VSS N_18 W=470n L=180.00n
MM2718 VSS WL<47> BL<2> VSS N_18 W=470n L=180.00n
MM2717 VSS WL<47> net4604 VSS N_18 W=470n L=180.00n
MM2716 VSS WL<47> net4608 VSS N_18 W=470n L=180.00n
MM2715 VSS WL<47> BL<4> VSS N_18 W=470n L=180.00n
MM2714 VSS WL<47> BL<6> VSS N_18 W=470n L=180.00n
MM2713 VSS WL<47> net4620 VSS N_18 W=470n L=180.00n
MM2712 VSS WL<47> net4624 VSS N_18 W=470n L=180.00n
MM2711 VSS WL<47> BL<8> VSS N_18 W=470n L=180.00n
MM2710 VSS WL<47> BL<10> VSS N_18 W=470n L=180.00n
MM2708 VSS WL<47> net4636 VSS N_18 W=470n L=180.00n
MM2707 VSS WL<47> net4640 VSS N_18 W=470n L=180.00n
MM2703 VSS WL<47> BL<14> VSS N_18 W=470n L=180.00n
MM2700 VSS WL<45> BL<14> VSS N_18 W=470n L=180.00n
MM2696 VSS WL<45> net4652 VSS N_18 W=470n L=180.00n
MM2695 VSS WL<45> net4656 VSS N_18 W=470n L=180.00n
MM2694 VSS WL<40> net4660 VSS N_18 W=470n L=180.00n
MM2692 VSS WL<45> BL<10> VSS N_18 W=470n L=180.00n
MM2691 VSS WL<45> BL<8> VSS N_18 W=470n L=180.00n
MM2690 VSS WL<45> net4672 VSS N_18 W=470n L=180.00n
MM2689 VSS WL<40> BL<13> VSS N_18 W=470n L=180.00n
MM2688 VSS WL<45> net4680 VSS N_18 W=470n L=180.00n
MM2687 VSS WL<40> BL<11> VSS N_18 W=470n L=180.00n
MM2686 VSS WL<45> BL<6> VSS N_18 W=470n L=180.00n
MM2685 VSS WL<45> BL<4> VSS N_18 W=470n L=180.00n
MM2684 VSS WL<45> net4696 VSS N_18 W=470n L=180.00n
MM2683 VSS WL<40> net4700 VSS N_18 W=470n L=180.00n
MM2682 VSS WL<45> net4704 VSS N_18 W=470n L=180.00n
MM2681 VSS WL<45> BL<2> VSS N_18 W=470n L=180.00n
MM2680 VSS WL<45> BL<0> VSS N_18 W=470n L=180.00n
MM2679 VSS WL<45> net4716 VSS N_18 W=470n L=180.00n
MM2671 VSS WL<43> BL<14> VSS N_18 W=470n L=180.00n
MM2670 VSS WL<45> BL<12> VSS N_18 W=470n L=180.00n
MM2666 VSS WL<45> net4728 VSS N_18 W=470n L=180.00n
MM2648 VSS WL<44> BL<15> VSS N_18 W=470n L=180.00n
MM2647 VSS WL<44> net4736 VSS N_18 W=470n L=180.00n
MM2646 VSS WL<44> net4740 VSS N_18 W=470n L=180.00n
MM2645 VSS WL<44> BL<13> VSS N_18 W=470n L=180.00n
MM2644 VSS WL<44> BL<11> VSS N_18 W=470n L=180.00n
MM2643 VSS WL<44> net4752 VSS N_18 W=470n L=180.00n
MM2642 VSS WL<44> net4756 VSS N_18 W=470n L=180.00n
MM2641 VSS WL<44> BL<9> VSS N_18 W=470n L=180.00n
MM2640 VSS WL<44> BL<7> VSS N_18 W=470n L=180.00n
MM2639 VSS WL<44> net4768 VSS N_18 W=470n L=180.00n
MM2638 VSS WL<44> net4772 VSS N_18 W=470n L=180.00n
MM2637 VSS WL<44> BL<5> VSS N_18 W=470n L=180.00n
MM2636 VSS WL<44> BL<3> VSS N_18 W=470n L=180.00n
MM2635 VSS WL<44> net4784 VSS N_18 W=470n L=180.00n
MM2634 VSS WL<44> BL<1> VSS N_18 W=470n L=180.00n
MM2633 VSS WL<44> net4792 VSS N_18 W=470n L=180.00n
MM2632 VSS WL<40> net4796 VSS N_18 W=470n L=180.00n
MM2631 VSS WL<40> BL<9> VSS N_18 W=470n L=180.00n
MM2629 VSS WL<40> BL<7> VSS N_18 W=470n L=180.00n
MM2628 VSS WL<40> net4808 VSS N_18 W=470n L=180.00n
MM2627 VSS WL<40> net4812 VSS N_18 W=470n L=180.00n
MM2626 VSS WL<40> BL<5> VSS N_18 W=470n L=180.00n
MM2625 VSS WL<41> BL<10> VSS N_18 W=470n L=180.00n
MM2624 VSS WL<41> BL<8> VSS N_18 W=470n L=180.00n
MM2623 VSS WL<41> net4828 VSS N_18 W=470n L=180.00n
MM2622 VSS WL<41> net4832 VSS N_18 W=470n L=180.00n
MM2621 VSS WL<41> BL<6> VSS N_18 W=470n L=180.00n
MM2620 VSS WL<41> BL<4> VSS N_18 W=470n L=180.00n
MM2619 VSS WL<41> net4844 VSS N_18 W=470n L=180.00n
MM2618 VSS WL<41> net4848 VSS N_18 W=470n L=180.00n
MM2617 VSS WL<41> BL<2> VSS N_18 W=470n L=180.00n
MM2616 VSS WL<41> BL<0> VSS N_18 W=470n L=180.00n
MM2615 VSS WL<43> net4860 VSS N_18 W=470n L=180.00n
MM2614 VSS WL<41> net4864 VSS N_18 W=470n L=180.00n
MM2613 VSS WL<43> BL<10> VSS N_18 W=470n L=180.00n
MM2611 VSS WL<40> BL<3> VSS N_18 W=470n L=180.00n
MM2609 VSS WL<43> net4876 VSS N_18 W=470n L=180.00n
MM2606 VSS WL<40> net4880 VSS N_18 W=470n L=180.00n
MM2597 VSS WL<41> BL<12> VSS N_18 W=470n L=180.00n
MM2593 VSS WL<41> net4888 VSS N_18 W=470n L=180.00n
MM2591 VSS WL<40> BL<1> VSS N_18 W=470n L=180.00n
MM2590 VSS WL<40> net4896 VSS N_18 W=470n L=180.00n
MM2589 VSS WL<56> net4900 VSS N_18 W=470n L=180.00n
MM2588 VSS WL<56> BL<1> VSS N_18 W=470n L=180.00n
MM2586 VSS WL<57> net4908 VSS N_18 W=470n L=180.00n
MM2582 VSS WL<57> BL<12> VSS N_18 W=470n L=180.00n
MM2573 VSS WL<56> net4916 VSS N_18 W=470n L=180.00n
MM2570 VSS WL<59> net4920 VSS N_18 W=470n L=180.00n
MM2568 VSS WL<56> BL<3> VSS N_18 W=470n L=180.00n
MM2566 VSS WL<59> BL<10> VSS N_18 W=470n L=180.00n
MM2565 VSS WL<57> net4932 VSS N_18 W=470n L=180.00n
MM2564 VSS WL<59> net4936 VSS N_18 W=470n L=180.00n
MM2563 VSS WL<57> BL<0> VSS N_18 W=470n L=180.00n
MM2562 VSS WL<57> BL<2> VSS N_18 W=470n L=180.00n
MM2561 VSS WL<57> net4948 VSS N_18 W=470n L=180.00n
MM2560 VSS WL<57> net4952 VSS N_18 W=470n L=180.00n
MM2559 VSS WL<57> BL<4> VSS N_18 W=470n L=180.00n
MM2558 VSS WL<57> BL<6> VSS N_18 W=470n L=180.00n
MM2557 VSS WL<57> net4964 VSS N_18 W=470n L=180.00n
MM2556 VSS WL<57> net4968 VSS N_18 W=470n L=180.00n
MM2555 VSS WL<57> BL<8> VSS N_18 W=470n L=180.00n
MM2554 VSS WL<57> BL<10> VSS N_18 W=470n L=180.00n
MM2553 VSS WL<56> BL<5> VSS N_18 W=470n L=180.00n
MM2552 VSS WL<56> net4984 VSS N_18 W=470n L=180.00n
MM2551 VSS WL<56> net4988 VSS N_18 W=470n L=180.00n
MM2550 VSS WL<56> BL<7> VSS N_18 W=470n L=180.00n
MM2548 VSS WL<56> BL<9> VSS N_18 W=470n L=180.00n
MM2547 VSS WL<56> net5000 VSS N_18 W=470n L=180.00n
MM2546 VSS WL<60> net5004 VSS N_18 W=470n L=180.00n
MM2545 VSS WL<60> BL<1> VSS N_18 W=470n L=180.00n
MM2544 VSS WL<60> net5012 VSS N_18 W=470n L=180.00n
MM2543 VSS WL<60> BL<3> VSS N_18 W=470n L=180.00n
MM2542 VSS WL<60> BL<5> VSS N_18 W=470n L=180.00n
MM2541 VSS WL<60> net5024 VSS N_18 W=470n L=180.00n
MM2540 VSS WL<60> net5028 VSS N_18 W=470n L=180.00n
MM2539 VSS WL<60> BL<7> VSS N_18 W=470n L=180.00n
MM2538 VSS WL<60> BL<9> VSS N_18 W=470n L=180.00n
MM2537 VSS WL<60> net5040 VSS N_18 W=470n L=180.00n
MM2536 VSS WL<60> net5044 VSS N_18 W=470n L=180.00n
MM2535 VSS WL<60> BL<11> VSS N_18 W=470n L=180.00n
MM2534 VSS WL<60> BL<13> VSS N_18 W=470n L=180.00n
MM2533 VSS WL<60> net5056 VSS N_18 W=470n L=180.00n
MM2532 VSS WL<60> net5060 VSS N_18 W=470n L=180.00n
MM2531 VSS WL<60> BL<15> VSS N_18 W=470n L=180.00n
MM2513 VSS WL<61> net5068 VSS N_18 W=470n L=180.00n
MM2509 VSS WL<61> BL<12> VSS N_18 W=470n L=180.00n
MM2508 VSS WL<59> BL<14> VSS N_18 W=470n L=180.00n
MM2500 VSS WL<61> net5080 VSS N_18 W=470n L=180.00n
MM2499 VSS WL<61> BL<0> VSS N_18 W=470n L=180.00n
MM2498 VSS WL<61> BL<2> VSS N_18 W=470n L=180.00n
MM2497 VSS WL<61> net5092 VSS N_18 W=470n L=180.00n
MM2496 VSS WL<56> net5096 VSS N_18 W=470n L=180.00n
MM3080 VSS WL<32> BL<3> VSS N_18 W=470n L=180.00n
MM3078 VSS WL<35> BL<10> VSS N_18 W=470n L=180.00n
MM3077 VSS WL<33> net5108 VSS N_18 W=470n L=180.00n
MM3076 VSS WL<35> net5112 VSS N_18 W=470n L=180.00n
MM3075 VSS WL<33> BL<0> VSS N_18 W=470n L=180.00n
MM3074 VSS WL<33> BL<2> VSS N_18 W=470n L=180.00n
MM3073 VSS WL<33> net5124 VSS N_18 W=470n L=180.00n
MM3072 VSS WL<33> net5128 VSS N_18 W=470n L=180.00n
MM3071 VSS WL<33> BL<4> VSS N_18 W=470n L=180.00n
MM3070 VSS WL<33> BL<6> VSS N_18 W=470n L=180.00n
MM3069 VSS WL<33> net5140 VSS N_18 W=470n L=180.00n
MM3068 VSS WL<33> net5144 VSS N_18 W=470n L=180.00n
MM3067 VSS WL<33> BL<8> VSS N_18 W=470n L=180.00n
MM3066 VSS WL<33> BL<10> VSS N_18 W=470n L=180.00n
MM3065 VSS WL<32> BL<5> VSS N_18 W=470n L=180.00n
MM3064 VSS WL<32> net5160 VSS N_18 W=470n L=180.00n
MM3063 VSS WL<32> net5164 VSS N_18 W=470n L=180.00n
MM3062 VSS WL<32> BL<7> VSS N_18 W=470n L=180.00n
MM3060 VSS WL<32> BL<9> VSS N_18 W=470n L=180.00n
MM3059 VSS WL<32> net5176 VSS N_18 W=470n L=180.00n
MM3058 VSS WL<36> net5180 VSS N_18 W=470n L=180.00n
MM3057 VSS WL<36> BL<1> VSS N_18 W=470n L=180.00n
MM3056 VSS WL<36> net5188 VSS N_18 W=470n L=180.00n
MM3055 VSS WL<36> BL<3> VSS N_18 W=470n L=180.00n
MM3054 VSS WL<36> BL<5> VSS N_18 W=470n L=180.00n
MM3053 VSS WL<36> net5200 VSS N_18 W=470n L=180.00n
MM3052 VSS WL<36> net5204 VSS N_18 W=470n L=180.00n
MM3051 VSS WL<36> BL<7> VSS N_18 W=470n L=180.00n
MM3050 VSS WL<36> BL<9> VSS N_18 W=470n L=180.00n
MM3049 VSS WL<36> net5216 VSS N_18 W=470n L=180.00n
MM3048 VSS WL<36> net5220 VSS N_18 W=470n L=180.00n
MM3047 VSS WL<36> BL<11> VSS N_18 W=470n L=180.00n
MM3046 VSS WL<36> BL<13> VSS N_18 W=470n L=180.00n
MM3045 VSS WL<36> net5232 VSS N_18 W=470n L=180.00n
MM3044 VSS WL<36> net5236 VSS N_18 W=470n L=180.00n
MM3043 VSS WL<36> BL<15> VSS N_18 W=470n L=180.00n
MM3025 VSS WL<37> net5244 VSS N_18 W=470n L=180.00n
MM3021 VSS WL<37> BL<12> VSS N_18 W=470n L=180.00n
MM3020 VSS WL<35> BL<14> VSS N_18 W=470n L=180.00n
MM3012 VSS WL<37> net5256 VSS N_18 W=470n L=180.00n
MM3011 VSS WL<37> BL<0> VSS N_18 W=470n L=180.00n
MM3010 VSS WL<37> BL<2> VSS N_18 W=470n L=180.00n
MM3009 VSS WL<37> net5268 VSS N_18 W=470n L=180.00n
MM3008 VSS WL<32> net5272 VSS N_18 W=470n L=180.00n
MM3007 VSS WL<37> net5276 VSS N_18 W=470n L=180.00n
MM3006 VSS WL<37> BL<4> VSS N_18 W=470n L=180.00n
MM3005 VSS WL<37> BL<6> VSS N_18 W=470n L=180.00n
MM3004 VSS WL<32> BL<11> VSS N_18 W=470n L=180.00n
MM3003 VSS WL<37> net5292 VSS N_18 W=470n L=180.00n
MM3002 VSS WL<32> BL<13> VSS N_18 W=470n L=180.00n
MM3001 VSS WL<37> net5300 VSS N_18 W=470n L=180.00n
MM3000 VSS WL<37> BL<8> VSS N_18 W=470n L=180.00n
MM2999 VSS WL<37> BL<10> VSS N_18 W=470n L=180.00n
MM2997 VSS WL<32> net5312 VSS N_18 W=470n L=180.00n
MM2996 VSS WL<37> net5316 VSS N_18 W=470n L=180.00n
MM2995 VSS WL<37> net5320 VSS N_18 W=470n L=180.00n
MM2991 VSS WL<37> BL<14> VSS N_18 W=470n L=180.00n
MM2988 VSS WL<39> BL<14> VSS N_18 W=470n L=180.00n
MM2984 VSS WL<39> net5332 VSS N_18 W=470n L=180.00n
MM2983 VSS WL<39> net5336 VSS N_18 W=470n L=180.00n
MM2981 VSS WL<39> BL<10> VSS N_18 W=470n L=180.00n
MM2980 VSS WL<39> BL<8> VSS N_18 W=470n L=180.00n
MM2979 VSS WL<39> net5348 VSS N_18 W=470n L=180.00n
MM2978 VSS WL<39> net5352 VSS N_18 W=470n L=180.00n
MM2977 VSS WL<39> BL<6> VSS N_18 W=470n L=180.00n
MM2976 VSS WL<39> BL<4> VSS N_18 W=470n L=180.00n
MM2975 VSS WL<39> net5364 VSS N_18 W=470n L=180.00n
MM2974 VSS WL<39> net5368 VSS N_18 W=470n L=180.00n
MM2973 VSS WL<39> BL<2> VSS N_18 W=470n L=180.00n
MM2972 VSS WL<39> BL<0> VSS N_18 W=470n L=180.00n
MM2971 VSS WL<39> net5380 VSS N_18 W=470n L=180.00n
MM2963 VSS WL<39> BL<12> VSS N_18 W=470n L=180.00n
MM2959 VSS WL<39> net5388 VSS N_18 W=470n L=180.00n
MM2948 VSS WL<33> net5392 VSS N_18 W=470n L=180.00n
MM2940 VSS WL<38> BL<15> VSS N_18 W=470n L=180.00n
MM2939 VSS WL<38> net5400 VSS N_18 W=470n L=180.00n
MM2938 VSS WL<38> net5404 VSS N_18 W=470n L=180.00n
MM2937 VSS WL<38> BL<13> VSS N_18 W=470n L=180.00n
MM2936 VSS WL<38> BL<11> VSS N_18 W=470n L=180.00n
MM2935 VSS WL<38> net5416 VSS N_18 W=470n L=180.00n
MM2934 VSS WL<38> net5420 VSS N_18 W=470n L=180.00n
MM2933 VSS WL<38> BL<9> VSS N_18 W=470n L=180.00n
MM2932 VSS WL<38> BL<7> VSS N_18 W=470n L=180.00n
MM2931 VSS WL<38> net5432 VSS N_18 W=470n L=180.00n
MM2930 VSS WL<38> net5436 VSS N_18 W=470n L=180.00n
MM2929 VSS WL<38> BL<5> VSS N_18 W=470n L=180.00n
MM2928 VSS WL<38> BL<3> VSS N_18 W=470n L=180.00n
MM2927 VSS WL<38> net5448 VSS N_18 W=470n L=180.00n
MM2926 VSS WL<38> BL<1> VSS N_18 W=470n L=180.00n
MM2925 VSS WL<38> net5456 VSS N_18 W=470n L=180.00n
MM2924 VSS WL<32> net5460 VSS N_18 W=470n L=180.00n
MM2923 VSS WL<32> BL<15> VSS N_18 W=470n L=180.00n
MM3101 VSS WL<32> net5468 VSS N_18 W=470n L=180.00n
MM3100 VSS WL<32> BL<1> VSS N_18 W=470n L=180.00n
MM3098 VSS WL<33> net5476 VSS N_18 W=470n L=180.00n
MM3094 VSS WL<33> BL<12> VSS N_18 W=470n L=180.00n
MM3085 VSS WL<32> net5484 VSS N_18 W=470n L=180.00n
MM3082 VSS WL<35> net5488 VSS N_18 W=470n L=180.00n
MM1329 VSS WL<11> BL<12> VSS N_18 W=470n L=180.00n
MM1333 VSS WL<11> net5496 VSS N_18 W=470n L=180.00n
MM1351 VSS WL<10> BL<15> VSS N_18 W=470n L=180.00n
MM1352 VSS WL<10> net5504 VSS N_18 W=470n L=180.00n
MM1353 VSS WL<10> net5508 VSS N_18 W=470n L=180.00n
MM1354 VSS WL<10> BL<13> VSS N_18 W=470n L=180.00n
MM1355 VSS WL<10> BL<11> VSS N_18 W=470n L=180.00n
MM1356 VSS WL<10> net5520 VSS N_18 W=470n L=180.00n
MM1357 VSS WL<10> net5524 VSS N_18 W=470n L=180.00n
MM1358 VSS WL<10> BL<9> VSS N_18 W=470n L=180.00n
MM1359 VSS WL<10> BL<7> VSS N_18 W=470n L=180.00n
MM1360 VSS WL<10> net5536 VSS N_18 W=470n L=180.00n
MM1361 VSS WL<10> net5540 VSS N_18 W=470n L=180.00n
MM1362 VSS WL<10> BL<5> VSS N_18 W=470n L=180.00n
MM1363 VSS WL<10> BL<3> VSS N_18 W=470n L=180.00n
MM1364 VSS WL<10> net5552 VSS N_18 W=470n L=180.00n
MM1365 VSS WL<10> BL<1> VSS N_18 W=470n L=180.00n
MM1366 VSS WL<10> net5560 VSS N_18 W=470n L=180.00n
MM1378 VSS WL<9> net5564 VSS N_18 W=470n L=180.00n
MM1387 VSS WL<8> BL<15> VSS N_18 W=470n L=180.00n
MM1388 VSS WL<8> net5572 VSS N_18 W=470n L=180.00n
MM1389 VSS WL<14> net5576 VSS N_18 W=470n L=180.00n
MM1390 VSS WL<14> BL<1> VSS N_18 W=470n L=180.00n
MM1391 VSS WL<14> net5584 VSS N_18 W=470n L=180.00n
MM1392 VSS WL<14> BL<3> VSS N_18 W=470n L=180.00n
MM1393 VSS WL<14> BL<5> VSS N_18 W=470n L=180.00n
MM1394 VSS WL<14> net5596 VSS N_18 W=470n L=180.00n
MM1395 VSS WL<14> net5600 VSS N_18 W=470n L=180.00n
MM1396 VSS WL<14> BL<7> VSS N_18 W=470n L=180.00n
MM1397 VSS WL<14> BL<9> VSS N_18 W=470n L=180.00n
MM1398 VSS WL<14> net5612 VSS N_18 W=470n L=180.00n
MM1399 VSS WL<14> net5616 VSS N_18 W=470n L=180.00n
MM1400 VSS WL<14> BL<11> VSS N_18 W=470n L=180.00n
MM1401 VSS WL<14> BL<13> VSS N_18 W=470n L=180.00n
MM1402 VSS WL<14> net5628 VSS N_18 W=470n L=180.00n
MM1403 VSS WL<14> net5632 VSS N_18 W=470n L=180.00n
MM1404 VSS WL<14> BL<15> VSS N_18 W=470n L=180.00n
MM1412 VSS WL<9> net5640 VSS N_18 W=470n L=180.00n
MM1423 VSS WL<15> net5644 VSS N_18 W=470n L=180.00n
MM1427 VSS WL<15> BL<12> VSS N_18 W=470n L=180.00n
MM1435 VSS WL<15> net5652 VSS N_18 W=470n L=180.00n
MM1436 VSS WL<15> BL<0> VSS N_18 W=470n L=180.00n
MM1437 VSS WL<15> BL<2> VSS N_18 W=470n L=180.00n
MM1438 VSS WL<15> net5664 VSS N_18 W=470n L=180.00n
MM1439 VSS WL<15> net5668 VSS N_18 W=470n L=180.00n
MM1440 VSS WL<15> BL<4> VSS N_18 W=470n L=180.00n
MM1441 VSS WL<15> BL<6> VSS N_18 W=470n L=180.00n
MM1442 VSS WL<15> net5680 VSS N_18 W=470n L=180.00n
MM1443 VSS WL<15> net5684 VSS N_18 W=470n L=180.00n
MM1444 VSS WL<15> BL<8> VSS N_18 W=470n L=180.00n
MM1445 VSS WL<15> BL<10> VSS N_18 W=470n L=180.00n
MM1447 VSS WL<15> net5696 VSS N_18 W=470n L=180.00n
MM1448 VSS WL<15> net5700 VSS N_18 W=470n L=180.00n
MM1452 VSS WL<15> BL<14> VSS N_18 W=470n L=180.00n
MM1455 VSS WL<13> BL<14> VSS N_18 W=470n L=180.00n
MM1104 VSS WL<1> BL<12> VSS N_18 W=470n L=180.00n
MM1459 VSS WL<13> net5716 VSS N_18 W=470n L=180.00n
MM1460 VSS WL<13> net5720 VSS N_18 W=470n L=180.00n
MM1461 VSS WL<8> net5724 VSS N_18 W=470n L=180.00n
MM1463 VSS WL<13> BL<10> VSS N_18 W=470n L=180.00n
MM1464 VSS WL<13> BL<8> VSS N_18 W=470n L=180.00n
MM1465 VSS WL<13> net5736 VSS N_18 W=470n L=180.00n
MM1466 VSS WL<8> BL<13> VSS N_18 W=470n L=180.00n
MM1467 VSS WL<13> net5744 VSS N_18 W=470n L=180.00n
MM1468 VSS WL<8> BL<11> VSS N_18 W=470n L=180.00n
MM1469 VSS WL<13> BL<6> VSS N_18 W=470n L=180.00n
MM1470 VSS WL<13> BL<4> VSS N_18 W=470n L=180.00n
MM1471 VSS WL<13> net5760 VSS N_18 W=470n L=180.00n
MM1472 VSS WL<8> net5764 VSS N_18 W=470n L=180.00n
MM1473 VSS WL<13> net5768 VSS N_18 W=470n L=180.00n
MM1474 VSS WL<13> BL<2> VSS N_18 W=470n L=180.00n
MM1475 VSS WL<13> BL<0> VSS N_18 W=470n L=180.00n
MM1476 VSS WL<13> net5780 VSS N_18 W=470n L=180.00n
MM1484 VSS WL<11> BL<14> VSS N_18 W=470n L=180.00n
MM1485 VSS WL<13> BL<12> VSS N_18 W=470n L=180.00n
MM1489 VSS WL<13> net5792 VSS N_18 W=470n L=180.00n
MM1102 VSS WL<1> net5796 VSS N_18 W=470n L=180.00n
MM1 VSS WL<0> BL<1> VSS N_18 W=470n L=180.00n
MM0 VSS WL<0> net5804 VSS N_18 W=470n L=180.00n
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    three_to8decoder_en
* View Name:    schematic
************************************************************************

.SUBCKT three_to8decoder_en A B C EN OUT0 OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 OUT7 
+ VDD VSS
*.PININFO A:I B:I C:I EN:I OUT0:O OUT1:O OUT2:O OUT3:O OUT4:O OUT5:O OUT6:O 
*.PININFO OUT7:O VDD:B VSS:B
XI7 A B C EN OUT7 VDD VSS / nand4
XI6 A B net0116 EN OUT6 VDD VSS / nand4
XI5 A net0105 C EN OUT5 VDD VSS / nand4
XI4 A net0105 net0116 EN OUT4 VDD VSS / nand4
XI3 net0158 B C EN OUT3 VDD VSS / nand4
XI2 net0158 B net0116 EN OUT2 VDD VSS / nand4
XI1 net0158 net0105 C EN OUT1 VDD VSS / nand4
XI0 net0158 net0105 net0116 EN OUT0 VDD VSS / nand4
XI11 B net0105 VDD VSS / inverter
XI10 C net0116 VDD VSS / inverter
XI8 A net0158 VDD VSS / inverter
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor A B OUT VDD VSS
*.PININFO A:I B:I OUT:O VDD:B VSS:B
MM5 OUT B VSS VSS N_18 W=500.0n L=180.00n m=1
MM4 OUT A VSS VSS N_18 W=500.0n L=180.00n m=1
MM10 net043 A VDD VDD P_18 W=500.0n L=180.00n m=3
MM0 OUT B net043 VDD P_18 W=500.0n L=180.00n m=3
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    six_to64decoder_en
* View Name:    schematic
************************************************************************

.SUBCKT six_to64decoder_en EN OUT<0> OUT<1> OUT<2> OUT<3> OUT<4> OUT<5> OUT<6> 
+ OUT<7> OUT<8> OUT<9> OUT<10> OUT<11> OUT<12> OUT<13> OUT<14> OUT<15> OUT<16> 
+ OUT<17> OUT<18> OUT<19> OUT<20> OUT<21> OUT<22> OUT<23> OUT<24> OUT<25> 
+ OUT<26> OUT<27> OUT<28> OUT<29> OUT<30> OUT<31> OUT<32> OUT<33> OUT<34> 
+ OUT<35> OUT<36> OUT<37> OUT<38> OUT<39> OUT<40> OUT<41> OUT<42> OUT<43> 
+ OUT<44> OUT<45> OUT<46> OUT<47> OUT<48> OUT<49> OUT<50> OUT<51> OUT<52> 
+ OUT<53> OUT<54> OUT<55> OUT<56> OUT<57> OUT<58> OUT<59> OUT<60> OUT<61> 
+ OUT<62> OUT<63> VDD VSS in0 in1 in2 in3 in4 in5
*.PININFO EN:I in0:I in1:I in2:I in3:I in4:I in5:I OUT<0>:O OUT<1>:O OUT<2>:O 
*.PININFO OUT<3>:O OUT<4>:O OUT<5>:O OUT<6>:O OUT<7>:O OUT<8>:O OUT<9>:O 
*.PININFO OUT<10>:O OUT<11>:O OUT<12>:O OUT<13>:O OUT<14>:O OUT<15>:O 
*.PININFO OUT<16>:O OUT<17>:O OUT<18>:O OUT<19>:O OUT<20>:O OUT<21>:O 
*.PININFO OUT<22>:O OUT<23>:O OUT<24>:O OUT<25>:O OUT<26>:O OUT<27>:O 
*.PININFO OUT<28>:O OUT<29>:O OUT<30>:O OUT<31>:O OUT<32>:O OUT<33>:O 
*.PININFO OUT<34>:O OUT<35>:O OUT<36>:O OUT<37>:O OUT<38>:O OUT<39>:O 
*.PININFO OUT<40>:O OUT<41>:O OUT<42>:O OUT<43>:O OUT<44>:O OUT<45>:O 
*.PININFO OUT<46>:O OUT<47>:O OUT<48>:O OUT<49>:O OUT<50>:O OUT<51>:O 
*.PININFO OUT<52>:O OUT<53>:O OUT<54>:O OUT<55>:O OUT<56>:O OUT<57>:O 
*.PININFO OUT<58>:O OUT<59>:O OUT<60>:O OUT<61>:O OUT<62>:O OUT<63>:O VDD:B 
*.PININFO VSS:B
XI1 in2 in1 in0 EN net11 net10 net9 net8 net7 net6 net5 net4 VDD VSS / 
+ three_to8decoder_en
XI0 in5 in4 in3 EN net24 net23 net22 net21 net20 net19 net18 net17 VDD VSS / 
+ three_to8decoder_en
XI146 net11 net18 OUT<48> VDD VSS / nor
XI145 net10 net18 OUT<49> VDD VSS / nor
XI144 net8 net18 OUT<51> VDD VSS / nor
XI143 net9 net18 OUT<50> VDD VSS / nor
XI142 net5 net18 OUT<54> VDD VSS / nor
XI141 net4 net18 OUT<55> VDD VSS / nor
XI140 net6 net18 OUT<53> VDD VSS / nor
XI139 net7 net18 OUT<52> VDD VSS / nor
XI138 net7 net17 OUT<60> VDD VSS / nor
XI137 net6 net17 OUT<61> VDD VSS / nor
XI136 net4 net17 OUT<63> VDD VSS / nor
XI135 net5 net17 OUT<62> VDD VSS / nor
XI134 net9 net17 OUT<58> VDD VSS / nor
XI121 net6 net20 OUT<37> VDD VSS / nor
XI120 net4 net20 OUT<39> VDD VSS / nor
XI119 net5 net20 OUT<38> VDD VSS / nor
XI118 net9 net20 OUT<34> VDD VSS / nor
XI117 net8 net20 OUT<35> VDD VSS / nor
XI116 net10 net20 OUT<33> VDD VSS / nor
XI115 net11 net20 OUT<32> VDD VSS / nor
XI84 net10 net24 OUT<1> VDD VSS / nor
XI85 net8 net24 OUT<3> VDD VSS / nor
XI86 net9 net24 OUT<2> VDD VSS / nor
XI87 net5 net24 OUT<6> VDD VSS / nor
XI88 net4 net24 OUT<7> VDD VSS / nor
XI89 net6 net24 OUT<5> VDD VSS / nor
XI90 net7 net24 OUT<4> VDD VSS / nor
XI91 net7 net23 OUT<12> VDD VSS / nor
XI92 net6 net23 OUT<13> VDD VSS / nor
XI93 net4 net23 OUT<15> VDD VSS / nor
XI94 net5 net23 OUT<14> VDD VSS / nor
XI95 net9 net23 OUT<10> VDD VSS / nor
XI96 net8 net23 OUT<11> VDD VSS / nor
XI97 net10 net23 OUT<9> VDD VSS / nor
XI98 net11 net23 OUT<8> VDD VSS / nor
XI132 net10 net17 OUT<57> VDD VSS / nor
XI131 net11 net17 OUT<56> VDD VSS / nor
XI130 net11 net19 OUT<40> VDD VSS / nor
XI129 net10 net19 OUT<41> VDD VSS / nor
XI128 net8 net19 OUT<43> VDD VSS / nor
XI127 net9 net19 OUT<42> VDD VSS / nor
XI126 net5 net19 OUT<46> VDD VSS / nor
XI125 net4 net19 OUT<47> VDD VSS / nor
XI124 net6 net19 OUT<45> VDD VSS / nor
XI123 net7 net19 OUT<44> VDD VSS / nor
XI122 net7 net20 OUT<36> VDD VSS / nor
XI99 net11 net21 OUT<24> VDD VSS / nor
XI100 net10 net21 OUT<25> VDD VSS / nor
XI101 net8 net21 OUT<27> VDD VSS / nor
XI102 net9 net21 OUT<26> VDD VSS / nor
XI103 net5 net21 OUT<30> VDD VSS / nor
XI104 net4 net21 OUT<31> VDD VSS / nor
XI105 net6 net21 OUT<29> VDD VSS / nor
XI106 net7 net21 OUT<28> VDD VSS / nor
XI107 net7 net22 OUT<20> VDD VSS / nor
XI108 net6 net22 OUT<21> VDD VSS / nor
XI109 net4 net22 OUT<23> VDD VSS / nor
XI110 net5 net22 OUT<22> VDD VSS / nor
XI111 net9 net22 OUT<18> VDD VSS / nor
XI112 net8 net22 OUT<19> VDD VSS / nor
XI113 net10 net22 OUT<17> VDD VSS / nor
XI114 net11 net22 OUT<16> VDD VSS / nor
XI2 net11 net24 OUT<0> VDD VSS / nor
XI133 net8 net17 OUT<59> VDD VSS / nor
.ENDS

************************************************************************
* Library Name: vlsi
* Cell Name:    Final_noSA
* View Name:    schematic
************************************************************************

.SUBCKT Final A<0> A<1> A<2> A<3> A<4> A<5> A<6> A<7> A<8> BL<0> BL<1> 
+ BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> 
+ BL<14> BL<15> CLK DL<0> DL<1> Dout<0> Dout<1> SAEN SO<0> SO<1> VDD VSS Vref 
+ WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> WL<6> WL<7> WL<8> WL<9> WL<10> WL<11> 
+ WL<12> WL<13> WL<14> WL<15> WL<16> WL<17> WL<18> WL<19> WL<20> WL<21> WL<22> 
+ WL<23> WL<24> WL<25> WL<26> WL<27> WL<28> WL<29> WL<30> WL<31> WL<32> WL<33> 
+ WL<34> WL<35> WL<36> WL<37> WL<38> WL<39> WL<40> WL<41> WL<42> WL<43> WL<44> 
+ WL<45> WL<46> WL<47> WL<48> WL<49> WL<50> WL<51> WL<52> WL<53> WL<54> WL<55> 
+ WL<56> WL<57> WL<58> WL<59> WL<60> WL<61> WL<62> WL<63> WLEN X_sel<0> 
+ X_sel<1> X_sel<2> X_sel<3> X_sel<4> X_sel<5> YOUT<0> YOUT<1> YOUT<2> YOUT<3> 
+ YOUT<4> YOUT<5> YOUT<6> YOUT<7> Y_sel<0> Y_sel<1> Y_sel<2>
*.PININFO A<0>:I A<1>:I A<2>:I A<3>:I A<4>:I A<5>:I A<6>:I A<7>:I A<8>:I CLK:I 
*.PININFO VDD:I VSS:I Vref:I Dout<0>:O Dout<1>:O SO<0>:O SO<1>:O BL<0>:B 
*.PININFO BL<1>:B BL<2>:B BL<3>:B BL<4>:B BL<5>:B BL<6>:B BL<7>:B BL<8>:B 
*.PININFO BL<9>:B BL<10>:B BL<11>:B BL<12>:B BL<13>:B BL<14>:B BL<15>:B 
*.PININFO DL<0>:B DL<1>:B SAEN:B WL<0>:B WL<1>:B WL<2>:B WL<3>:B WL<4>:B 
*.PININFO WL<5>:B WL<6>:B WL<7>:B WL<8>:B WL<9>:B WL<10>:B WL<11>:B WL<12>:B 
*.PININFO WL<13>:B WL<14>:B WL<15>:B WL<16>:B WL<17>:B WL<18>:B WL<19>:B 
*.PININFO WL<20>:B WL<21>:B WL<22>:B WL<23>:B WL<24>:B WL<25>:B WL<26>:B 
*.PININFO WL<27>:B WL<28>:B WL<29>:B WL<30>:B WL<31>:B WL<32>:B WL<33>:B 
*.PININFO WL<34>:B WL<35>:B WL<36>:B WL<37>:B WL<38>:B WL<39>:B WL<40>:B 
*.PININFO WL<41>:B WL<42>:B WL<43>:B WL<44>:B WL<45>:B WL<46>:B WL<47>:B 
*.PININFO WL<48>:B WL<49>:B WL<50>:B WL<51>:B WL<52>:B WL<53>:B WL<54>:B 
*.PININFO WL<55>:B WL<56>:B WL<57>:B WL<58>:B WL<59>:B WL<60>:B WL<61>:B 
*.PININFO WL<62>:B WL<63>:B WLEN:B X_sel<0>:B X_sel<1>:B X_sel<2>:B X_sel<3>:B 
*.PININFO X_sel<4>:B X_sel<5>:B YOUT<0>:B YOUT<1>:B YOUT<2>:B YOUT<3>:B 
*.PININFO YOUT<4>:B YOUT<5>:B YOUT<6>:B YOUT<7>:B Y_sel<0>:B Y_sel<1>:B 
*.PININFO Y_sel<2>:B
XI29 A<0> A<1> A<2> A<3> A<4> A<5> A<6> A<7> A<8> CLK SAEN VDD VSS WLEN 
+ X_sel<0> X_sel<1> X_sel<2> X_sel<3> X_sel<4> X_sel<5> Y_sel<0> Y_sel<1> 
+ Y_sel<2> / timing_control2
XI27 SAEN DL<0> Vref SO<0> Dout<0> VDD VSS / SA_Final
XI28 SAEN DL<1> Vref SO<1> Dout<1> VDD VSS / SA_Final
XI26 Y_sel<0> Y_sel<1> Y_sel<2> VDD YOUT<0> YOUT<1> YOUT<2> YOUT<3> YOUT<4> 
+ YOUT<5> YOUT<6> YOUT<7> VDD VSS / to8decoder_en
XI17 BL<8> BL<9> BL<10> BL<11> BL<12> BL<13> BL<14> BL<15> DL<1> VDD VSS 
+ YOUT<0> YOUT<1> YOUT<2> YOUT<3> YOUT<4> YOUT<5> YOUT<6> YOUT<7> / YMUX
XI16 BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> DL<0> VDD VSS YOUT<0> 
+ YOUT<1> YOUT<2> YOUT<3> YOUT<4> YOUT<5> YOUT<6> YOUT<7> / YMUX
XI13 BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> 
+ BL<12> BL<13> BL<14> BL<15> VDD CLK / precharge
XI10 BL<0> BL<1> BL<2> BL<3> BL<4> BL<5> BL<6> BL<7> BL<8> BL<9> BL<10> BL<11> 
+ BL<12> BL<13> BL<14> BL<15> VSS WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> WL<6> 
+ WL<7> WL<8> WL<9> WL<10> WL<11> WL<12> WL<13> WL<14> WL<15> WL<16> WL<17> 
+ WL<18> WL<19> WL<20> WL<21> WL<22> WL<23> WL<24> WL<25> WL<26> WL<27> WL<28> 
+ WL<29> WL<30> WL<31> WL<32> WL<33> WL<34> WL<35> WL<36> WL<37> WL<38> WL<39> 
+ WL<40> WL<41> WL<42> WL<43> WL<44> WL<45> WL<46> WL<47> WL<48> WL<49> WL<50> 
+ WL<51> WL<52> WL<53> WL<54> WL<55> WL<56> WL<57> WL<58> WL<59> WL<60> WL<61> 
+ WL<62> WL<63> / ROM
XI9 WLEN WL<0> WL<1> WL<2> WL<3> WL<4> WL<5> WL<6> WL<7> WL<8> WL<9> WL<10> 
+ WL<11> WL<12> WL<13> WL<14> WL<15> WL<16> WL<17> WL<18> WL<19> WL<20> WL<21> 
+ WL<22> WL<23> WL<24> WL<25> WL<26> WL<27> WL<28> WL<29> WL<30> WL<31> WL<32> 
+ WL<33> WL<34> WL<35> WL<36> WL<37> WL<38> WL<39> WL<40> WL<41> WL<42> WL<43> 
+ WL<44> WL<45> WL<46> WL<47> WL<48> WL<49> WL<50> WL<51> WL<52> WL<53> WL<54> 
+ WL<55> WL<56> WL<57> WL<58> WL<59> WL<60> WL<61> WL<62> WL<63> VDD VSS 
+ X_sel<0> X_sel<1> X_sel<2> X_sel<3> X_sel<4> X_sel<5> / six_to64decoder_en
.ENDS

