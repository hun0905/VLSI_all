* SPICE NETLIST
***************************************

.SUBCKT RM1 A B
.ENDS
***************************************
.SUBCKT RM2 A B
.ENDS
***************************************
.SUBCKT RM3 A B
.ENDS
***************************************
.SUBCKT RM4 A B
.ENDS
***************************************
.SUBCKT RM5 A B
.ENDS
***************************************
.SUBCKT RM6 A B
.ENDS
***************************************
.SUBCKT DN A B
.ENDS
***************************************
.SUBCKT DP A B
.ENDS
***************************************
.SUBCKT L_SLCR20K_RF POS NEG SUB
.ENDS
***************************************
.SUBCKT PAD_RF POS NEG
.ENDS
***************************************
.SUBCKT nmos_small
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_small
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT hw2_part1_2 VSS A B VDD C OUT
** N=8 EP=6 IP=720 FDC=39
M0 OUT A 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=-1070 $Y=2660 $D=0
M1 4 A OUT VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=-380 $Y=2660 $D=0
M2 OUT A 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=310 $Y=2660 $D=0
M3 4 A OUT VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=1000 $Y=2660 $D=0
M4 OUT A 4 VSS N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=1690 $Y=2660 $D=0
M5 VSS B 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=3250 $Y=2660 $D=0
M6 4 B VSS VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=3940 $Y=2660 $D=0
M7 VSS B 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=4630 $Y=2660 $D=0
M8 4 B VSS VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=5320 $Y=2660 $D=0
M9 VSS B 4 VSS N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=6010 $Y=2660 $D=0
M10 VSS C OUT VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=7570 $Y=2660 $D=0
M11 OUT C VSS VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=8260 $Y=2660 $D=0
M12 VSS C OUT VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=8950 $Y=2660 $D=0
M13 OUT C VSS VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=9640 $Y=2660 $D=0
M14 VSS C OUT VSS N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=10330 $Y=2660 $D=0
M15 8 A VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06 $X=-8275 $Y=9582 $D=1
M16 VDD A 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-7585 $Y=9582 $D=1
M17 8 A VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-6895 $Y=9582 $D=1
M18 VDD A 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-6205 $Y=9582 $D=1
M19 8 A VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-5515 $Y=9582 $D=1
M20 VDD A 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-4825 $Y=9582 $D=1
M21 8 A VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-4135 $Y=9582 $D=1
M22 VDD A 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-3445 $Y=9582 $D=1
M23 8 A VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-2755 $Y=9582 $D=1
M24 VDD A 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-2065 $Y=9582 $D=1
M25 8 A VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=-1375 $Y=9582 $D=1
M26 VDD A 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07 $X=-685 $Y=9582 $D=1
M27 8 B VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06 $X=1475 $Y=9584 $D=1
M28 VDD B 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=2165 $Y=9584 $D=1
M29 8 B VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=2855 $Y=9584 $D=1
M30 VDD B 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=3545 $Y=9584 $D=1
M31 8 B VDD VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=4235 $Y=9584 $D=1
M32 VDD B 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07 $X=4925 $Y=9584 $D=1
M33 OUT C 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=1.225e-12 PD=5.1e-07 PS=3.48e-06 $X=7085 $Y=9582 $D=1
M34 8 C OUT VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=7775 $Y=9582 $D=1
M35 OUT C 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=8465 $Y=9582 $D=1
M36 8 C OUT VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=9155 $Y=9582 $D=1
M37 OUT C 8 VDD P_18 L=1.8e-07 W=2.5e-06 AD=6.375e-13 AS=6.375e-13 PD=5.1e-07 PS=5.1e-07 $X=9845 $Y=9582 $D=1
M38 8 C OUT VDD P_18 L=1.8e-07 W=2.5e-06 AD=1.225e-12 AS=6.375e-13 PD=3.48e-06 PS=5.1e-07 $X=10535 $Y=9582 $D=1
.ENDS
***************************************
