* SPICE NETLIST
***************************************

*.CALIBRE ABORT_INFO SOFTCHK
.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT nmos_small
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_small
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT hw2_part1_1 C B VDD A VSS OUT
** N=10 EP=6 IP=336 FDC=24
M0 VSS C 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=1690 $Y=-1235 $D=0
M1 4 C VSS VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=2380 $Y=-1235 $D=0
M2 VSS C 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=3070 $Y=-1235 $D=0
M3 4 C VSS VSS N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=3760 $Y=-1235 $D=0
M4 1 B 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=5320 $Y=-1235 $D=0
M5 4 B 1 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=6010 $Y=-1235 $D=0
M6 1 B 4 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=6700 $Y=-1235 $D=0
M7 4 B 1 VSS N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=7390 $Y=-1235 $D=0
M8 1 A OUT VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07 PS=2.98e-06 $X=10350 $Y=-1335 $D=0
M9 OUT A 1 VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=11040 $Y=-1335 $D=0
M10 1 A OUT VSS N_18 L=1.8e-07 W=2e-06 AD=5.1e-13 AS=5.1e-13 PD=5.1e-07 PS=5.1e-07 $X=11730 $Y=-1335 $D=0
M11 OUT A 1 VSS N_18 L=1.8e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06 PS=5.1e-07 $X=12420 $Y=-1335 $D=0
M12 OUT C VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=910 $Y=5220 $D=1
M13 OUT B VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06 $X=3070 $Y=5220 $D=1
M14 OUT A VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07 PS=2.48e-06 $X=5230 $Y=5220 $D=1
M15 VDD A OUT VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=5920 $Y=5220 $D=1
M16 OUT A VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=6610 $Y=5220 $D=1
M17 VDD A OUT VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=7300 $Y=5220 $D=1
M18 OUT A VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=7990 $Y=5220 $D=1
M19 VDD A OUT VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=8680 $Y=5220 $D=1
M20 OUT A VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=9370 $Y=5220 $D=1
M21 VDD A OUT VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=10060 $Y=5220 $D=1
M22 OUT A VDD VDD P_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=3.825e-13 PD=5.1e-07 PS=5.1e-07 $X=10750 $Y=5220 $D=1
M23 VDD A OUT VDD P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06 PS=5.1e-07 $X=11440 $Y=5220 $D=1
*.CALIBRE WARNING SCONNECT SCONNECT conflict(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
